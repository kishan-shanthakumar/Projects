module bintobcd(
input [3:0] i,
output reg [13:0] op);

always @(*)
begin
	case (i)
	4'b0000 : op = 14'b00000000111111;
	4'b0001 : op = 14'b00000000000110;
	4'b0010 : op = 14'b00000001011011;
	4'b0011 : op = 14'b00000001001111;
	4'b0100 : op = 14'b00000001100110;
	4'b0101 : op = 14'b00000001101101;
	4'b0110 : op = 14'b00000001111101;
	4'b0111 : op = 14'b00000000000111;
	4'b1000 : op = 14'b00000001111111;
	4'b1001 : op = 14'b00000001101111;
	4'b1010 : op = 14'b00001100111111;
	4'b1011 : op = 14'b00001100000110;
	4'b1100 : op = 14'b00001101011011;
	4'b1101 : op = 14'b00001101001111;
	4'b1110 : op = 14'b00001101100110;
	4'b1111 : op = 14'b00001101101101;
	endcase
	op = op ^ 14'b11111111111111;
end

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.08.2021 19:38:20
// Design Name: 
// Module Name: ham80_64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ham80_64(inp,outp);
input [79:0] inp;
output reg [15:0] outp;

reg [15:0] hmat[79:0];
reg [15:0] o;

integer temp;
integer i;
integer j;

initial begin
hmat[0] = 16'b0110000010010111;
hmat[1] = 16'b1111011010111101;
hmat[2] = 16'b1011110110101000;
hmat[3] = 16'b0101111011010100;
hmat[4] = 16'b0010111101101010;
hmat[5] = 16'b0001011110110101;
hmat[6] = 16'b1100110100101100;
hmat[7] = 16'b0110011010010110;
hmat[8] = 16'b0011001101001011;
hmat[9] = 16'b1101111101010011;
hmat[10] = 16'b1010100101011111;
hmat[11] = 16'b1001001001011001;
hmat[12] = 16'b1000111111011010;
hmat[13] = 16'b0100011111101101;
hmat[14] = 16'b1110010100000000;
hmat[15] = 16'b0111001010000000;
hmat[16] = 16'b0011100101000000;
hmat[17] = 16'b0001110010100000;
hmat[18] = 16'b0000111001010000;
hmat[19] = 16'b0000011100101000;
hmat[20] = 16'b0000001110010100;
hmat[21] = 16'b0000000111001010;
hmat[22] = 16'b0000000011100101;
hmat[23] = 16'b1100011010000100;
hmat[24] = 16'b0110001101000010;
hmat[25] = 16'b0011000110100001;
hmat[26] = 16'b1101111000100110;
hmat[27] = 16'b0110111100010011;
hmat[28] = 16'b1111000101111111;
hmat[29] = 16'b1011111001001001;
hmat[30] = 16'b1001100111010010;
hmat[31] = 16'b0100110011101001;
hmat[32] = 16'b1110000010000010;
hmat[33] = 16'b0111000001000001;
hmat[34] = 16'b1111111011010110;
hmat[35] = 16'b0111111101101011;
hmat[36] = 16'b1111100101000011;
hmat[37] = 16'b1011101001010111;
hmat[38] = 16'b1001101111011101;
hmat[39] = 16'b1000101100011000;
hmat[40] = 16'b0100010110001100;
hmat[41] = 16'b0010001011000110;
hmat[42] = 16'b0001000101100011;
hmat[43] = 16'b1100111001000111;
hmat[44] = 16'b1010000111010101;
hmat[45] = 16'b1001011000011100;
hmat[46] = 16'b0100101100001110;
hmat[47] = 16'b0010010110000111;
hmat[48] = 16'b1101010000110101;
hmat[49] = 16'b1010110011101100;
hmat[50] = 16'b0101011001110110;
hmat[51] = 16'b0010101100111011;
hmat[52] = 16'b1101001101101011;
hmat[53] = 16'b1010111101000011;
hmat[54] = 16'b1001000101010111;
hmat[55] = 16'b1000111001011101;
hmat[56] = 16'b1000000111011000;
hmat[57] = 16'b0100000011101100;
hmat[58] = 16'b0010000001110110;
hmat[59] = 16'b0001000000111011;
hmat[60] = 16'b1100111011101011;
hmat[61] = 16'b1010000110000011;
hmat[62] = 16'b1001011000110111;
hmat[63] = 16'b1000110111101101;
hmat[64] = 16'b1000000000000000;
hmat[65] = 16'b0100000000000000;
hmat[66] = 16'b0010000000000000;
hmat[67] = 16'b0001000000000000;
hmat[68] = 16'b0000100000000000;
hmat[69] = 16'b0000010000000000;
hmat[70] = 16'b0000001000000000;
hmat[71] = 16'b0000000100000000;
hmat[72] = 16'b0000000010000000;
hmat[73] = 16'b0000000001000000;
hmat[74] = 16'b0000000000100000;
hmat[75] = 16'b0000000000010000;
hmat[76] = 16'b0000000000001000;
hmat[77] = 16'b0000000000000100;
hmat[78] = 16'b0000000000000010;
hmat[79] = 16'b0000000000000001;
end

always @(*)
begin
    for(i = 0; i < 16; i = i + 1)
    begin
        temp = 0;
        for(j = 0; j < 80; j = j + 1)
        begin
            temp = temp ^ (hmat[j][15-i] & inp[79-j]);
        end
        o[15-i] = temp;
    end
    outp = o;
end

endmodule

module sub(input [7:0] sub_a,sub_b,
			output [7:0] diff);

assign diff = sub_a - sub_b;

endmodule
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.08.2021 17:46:19
// Design Name: 
// Module Name: ham80_64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module ham80_64e(inp, outp);
input [63:0] inp;
output reg [79:0] outp;

reg [79:0] gen[63:0];
reg [79:0] o;

integer temp;
integer i;
integer j;

initial begin
gen[0]  = 80'b10000000000000000000000000000000000000000000000000000000000000000110000010010111;
gen[1]  = 80'b01000000000000000000000000000000000000000000000000000000000000001111011010111101;
gen[2]  = 80'b00100000000000000000000000000000000000000000000000000000000000001011110110101000;
gen[3]  = 80'b00010000000000000000000000000000000000000000000000000000000000000101111011010100;
gen[4]  = 80'b00001000000000000000000000000000000000000000000000000000000000000010111101101010;
gen[5]  = 80'b00000100000000000000000000000000000000000000000000000000000000000001011110110101;
gen[6]  = 80'b00000010000000000000000000000000000000000000000000000000000000001100110100101100;
gen[7]  = 80'b00000001000000000000000000000000000000000000000000000000000000000110011010010110;
gen[8]  = 80'b00000000100000000000000000000000000000000000000000000000000000000011001101001011;
gen[9]  = 80'b00000000010000000000000000000000000000000000000000000000000000001101111101010011;
gen[10] = 80'b00000000001000000000000000000000000000000000000000000000000000001010100101011111;
gen[11] = 80'b00000000000100000000000000000000000000000000000000000000000000001001001001011001;
gen[12] = 80'b00000000000010000000000000000000000000000000000000000000000000001000111111011010;
gen[13] = 80'b00000000000001000000000000000000000000000000000000000000000000000100011111101101;
gen[14] = 80'b00000000000000100000000000000000000000000000000000000000000000001110010100000000;
gen[15] = 80'b00000000000000010000000000000000000000000000000000000000000000000111001010000000;
gen[16] = 80'b00000000000000001000000000000000000000000000000000000000000000000011100101000000;
gen[17] = 80'b00000000000000000100000000000000000000000000000000000000000000000001110010100000;
gen[18] = 80'b00000000000000000010000000000000000000000000000000000000000000000000111001010000;
gen[19] = 80'b00000000000000000001000000000000000000000000000000000000000000000000011100101000;
gen[20] = 80'b00000000000000000000100000000000000000000000000000000000000000000000001110010100;
gen[21] = 80'b00000000000000000000010000000000000000000000000000000000000000000000000111001010;
gen[22] = 80'b00000000000000000000001000000000000000000000000000000000000000000000000011100101;
gen[23] = 80'b00000000000000000000000100000000000000000000000000000000000000001100011010000100;
gen[24] = 80'b00000000000000000000000010000000000000000000000000000000000000000110001101000010;
gen[25] = 80'b00000000000000000000000001000000000000000000000000000000000000000011000110100001;
gen[26] = 80'b00000000000000000000000000100000000000000000000000000000000000001101111000100110;
gen[27] = 80'b00000000000000000000000000010000000000000000000000000000000000000110111100010011;
gen[28] = 80'b00000000000000000000000000001000000000000000000000000000000000001111000101111111;
gen[29] = 80'b00000000000000000000000000000100000000000000000000000000000000001011111001001001;
gen[30] = 80'b00000000000000000000000000000010000000000000000000000000000000001001100111010010;
gen[31] = 80'b00000000000000000000000000000001000000000000000000000000000000000100110011101001;
gen[32] = 80'b00000000000000000000000000000000100000000000000000000000000000001110000010000010;
gen[33] = 80'b00000000000000000000000000000000010000000000000000000000000000000111000001000001;
gen[34] = 80'b00000000000000000000000000000000001000000000000000000000000000001111111011010110;
gen[35] = 80'b00000000000000000000000000000000000100000000000000000000000000000111111101101011;
gen[36] = 80'b00000000000000000000000000000000000010000000000000000000000000001111100101000011;
gen[37] = 80'b00000000000000000000000000000000000001000000000000000000000000001011101001010111;
gen[38] = 80'b00000000000000000000000000000000000000100000000000000000000000001001101111011101;
gen[39] = 80'b00000000000000000000000000000000000000010000000000000000000000001000101100011000;
gen[40] = 80'b00000000000000000000000000000000000000001000000000000000000000000100010110001100;
gen[41] = 80'b00000000000000000000000000000000000000000100000000000000000000000010001011000110;
gen[42] = 80'b00000000000000000000000000000000000000000010000000000000000000000001000101100011;
gen[43] = 80'b00000000000000000000000000000000000000000001000000000000000000001100111001000111;
gen[44] = 80'b00000000000000000000000000000000000000000000100000000000000000001010000111010101;
gen[45] = 80'b00000000000000000000000000000000000000000000010000000000000000001001011000011100;
gen[46] = 80'b00000000000000000000000000000000000000000000001000000000000000000100101100001110;
gen[47] = 80'b00000000000000000000000000000000000000000000000100000000000000000010010110000111;
gen[48] = 80'b00000000000000000000000000000000000000000000000010000000000000001101010000110101;
gen[49] = 80'b00000000000000000000000000000000000000000000000001000000000000001010110011101100;
gen[50] = 80'b00000000000000000000000000000000000000000000000000100000000000000101011001110110;
gen[51] = 80'b00000000000000000000000000000000000000000000000000010000000000000010101100111011;
gen[52] = 80'b00000000000000000000000000000000000000000000000000001000000000001101001101101011;
gen[53] = 80'b00000000000000000000000000000000000000000000000000000100000000001010111101000011;
gen[54] = 80'b00000000000000000000000000000000000000000000000000000010000000001001000101010111;
gen[55] = 80'b00000000000000000000000000000000000000000000000000000001000000001000111001011101;
gen[56] = 80'b00000000000000000000000000000000000000000000000000000000100000001000000111011000;
gen[57] = 80'b00000000000000000000000000000000000000000000000000000000010000000100000011101100;
gen[58] = 80'b00000000000000000000000000000000000000000000000000000000001000000010000001110110;
gen[59] = 80'b00000000000000000000000000000000000000000000000000000000000100000001000000111011;
gen[60] = 80'b00000000000000000000000000000000000000000000000000000000000010001100111011101011;
gen[61] = 80'b00000000000000000000000000000000000000000000000000000000000001001010000110000011;
gen[62] = 80'b00000000000000000000000000000000000000000000000000000000000000101001011000110111;
gen[63] = 80'b00000000000000000000000000000000000000000000000000000000000000011000110111101101;
end

always @(*)
begin
    for(i = 0; i < 80; i = i + 1)
    begin
        temp = 0;
        for(j = 0; j < 64; j = j + 1)
        begin
            temp = temp ^ (gen[j][79-i] & inp[63-j]);
        end
        o[79-i] = temp;
    end
    outp = o;
end

endmodule

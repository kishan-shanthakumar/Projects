module spi();
endmodule

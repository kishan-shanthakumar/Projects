module usb2();
endmodule

module riscv_core();
output [31:0] addr;
input [31:0] dout;
output [31:0] din;

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07.09.2021 13:42:18
// Design Name: 
// Module Name: ham_4be
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ham_4be(
input [79:0] code,
input [15:0] syndrome,
output reg [63:0] dataout,
output reg ec
);

reg [79:0] data;

always @(*)
begin    
    case(syndrome)
        16'b0000000000000000:begin data = code; ec = 1; end
        16'b0000000000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0000000000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0000000000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0000000000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0000000000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0000000000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0000000001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0000000010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0000000100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0000001000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0000010000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0000100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0001000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0010000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0100000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1000000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1000110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1001011000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1010000110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1100111011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0001000000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0010000001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0100000011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1000000111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1000111001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1001000101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1010111101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1101001101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0010101100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0101011001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1010110011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1101010000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0010010110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0100101100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1001011000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1010000111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1100111001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0001000101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0010001011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0100010110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1000101100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1001101111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1011101001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000000000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000111; ec = 1; end
        16'b0000000000001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001110; ec = 1; end
        16'b0000000000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000011100; ec = 1; end
        16'b0000000000111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000111000; ec = 1; end
        16'b0000000001110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001110000; ec = 1; end
        16'b0000000011100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000011100000; ec = 1; end
        16'b0000000111000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000111000000; ec = 1; end
        16'b0000001110000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001110000000; ec = 1; end
        16'b0000011100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000011100000000; ec = 1; end
        16'b0000111000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000111000000000; ec = 1; end
        16'b0001110000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001110000000000; ec = 1; end
        16'b0011100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000011100000000000; ec = 1; end
        16'b0111000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000111000000000000; ec = 1; end
        16'b1110000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001110000000000000; ec = 1; end
        16'b0100110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000011100000000000000; ec = 1; end
        16'b1001101111011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000111000000000000000; ec = 1; end
        16'b1011101001011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001110000000000000000; ec = 1; end
        16'b1111100101011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000011100000000000000000; ec = 1; end
        16'b0111111101010011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000111000000000000000000; ec = 1; end
        16'b1111111010100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001110000000000000000000; ec = 1; end
        16'b0111000010100001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000011100000000000000000000; ec = 1; end
        16'b1110000101000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000111000000000000000000000; ec = 1; end
        16'b0100111101101001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001110000000000000000000000; ec = 1; end
        16'b1001111011010010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000011100000000000000000000000; ec = 1; end
        16'b1011000001001001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000111000000000000000000000000; ec = 1; end
        16'b1110110101111111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001110000000000000000000000000; ec = 1; end
        16'b0101011100010011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000011100000000000000000000000000; ec = 1; end
        16'b1010111000100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000111000000000000000000000000000; ec = 1; end
        16'b1101000110100001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001110000000000000000000000000000; ec = 1; end
        16'b0010111010101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000011100000000000000000000000000000; ec = 1; end
        16'b0101110101011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000111000000000000000000000000000000; ec = 1; end
        16'b1011101010111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000001110000000000000000000000000000000; ec = 1; end
        16'b1111100010010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000011100000000000000000000000000000000; ec = 1; end
        16'b0111110011000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000111000000000000000000000000000000000; ec = 1; end
        16'b1111100110001110:begin data = code ^ 80'b00000000000000000000000000000000000000000001110000000000000000000000000000000000; ec = 1; end
        16'b0111111011110001:begin data = code ^ 80'b00000000000000000000000000000000000000000011100000000000000000000000000000000000; ec = 1; end
        16'b1111110111100010:begin data = code ^ 80'b00000000000000000000000000000000000000000111000000000000000000000000000000000000; ec = 1; end
        16'b0111011000101001:begin data = code ^ 80'b00000000000000000000000000000000000000001110000000000000000000000000000000000000; ec = 1; end
        16'b1110110001010010:begin data = code ^ 80'b00000000000000000000000000000000000000011100000000000000000000000000000000000000; ec = 1; end
        16'b0101010101001001:begin data = code ^ 80'b00000000000000000000000000000000000000111000000000000000000000000000000000000000; ec = 1; end
        16'b1010101010010010:begin data = code ^ 80'b00000000000000000000000000000000000001110000000000000000000000000000000000000000; ec = 1; end
        16'b1101100011001001:begin data = code ^ 80'b00000000000000000000000000000000000011100000000000000000000000000000000000000000; ec = 1; end
        16'b0011110001111111:begin data = code ^ 80'b00000000000000000000000000000000000111000000000000000000000000000000000000000000; ec = 1; end
        16'b0111100011111110:begin data = code ^ 80'b00000000000000000000000000000000001110000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000111111100:begin data = code ^ 80'b00000000000000000000000000000000011100000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111000010101:begin data = code ^ 80'b00000000000000000000000000000000111000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101110000101010:begin data = code ^ 80'b00000000000000000000000000000001110000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011010110111001:begin data = code ^ 80'b00000000000000000000000000000011100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110101101110010:begin data = code ^ 80'b00000000000000000000000000000111000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101011011100100:begin data = code ^ 80'b00000000000000000000000000001110000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000000100101:begin data = code ^ 80'b00000000000000000000000000011100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100000001001010:begin data = code ^ 80'b00000000000000000000000000111000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000010010100:begin data = code ^ 80'b00000000000000000000000001110000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000110011000101:begin data = code ^ 80'b00000000000000000000000011100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001010001100111:begin data = code ^ 80'b00000000000000000000000111000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010010100100011:begin data = code ^ 80'b00000000000000000000001110000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011110101011:begin data = code ^ 80'b00000000000000000000011100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001010111011:begin data = code ^ 80'b00000000000000000000111000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000010101110110:begin data = code ^ 80'b00000000000000000001110000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101011101100:begin data = code ^ 80'b00000000000000000011100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001010111011000:begin data = code ^ 80'b00000000000000000111000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010101110110000:begin data = code ^ 80'b00000000000000001110000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101011101100000:begin data = code ^ 80'b00000000000000011100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111011000000:begin data = code ^ 80'b00000000000000111000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000001101101:begin data = code ^ 80'b00000000000001110000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110100110111:begin data = code ^ 80'b00000000000011100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101101001101110:begin data = code ^ 80'b00000000000111000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011010011011100:begin data = code ^ 80'b00000000001110000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010001010101:begin data = code ^ 80'b00000000011100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100010101000111:begin data = code ^ 80'b00000000111000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101010001110:begin data = code ^ 80'b00000001110000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100011110001:begin data = code ^ 80'b00000011100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110000001111:begin data = code ^ 80'b00000111000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111010111110011:begin data = code ^ 80'b00001110000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011000001011:begin data = code ^ 80'b00011100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110000010110:begin data = code ^ 80'b00111000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001010111000001:begin data = code ^ 80'b01110000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010101110000010:begin data = code ^ 80'b11100000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000000001011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001011; ec = 1; end
        16'b0000000000010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010110; ec = 1; end
        16'b0000000000101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000101100; ec = 1; end
        16'b0000000001011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001011000; ec = 1; end
        16'b0000000010110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010110000; ec = 1; end
        16'b0000000101100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000101100000; ec = 1; end
        16'b0000001011000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001011000000; ec = 1; end
        16'b0000010110000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010110000000; ec = 1; end
        16'b0000101100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000101100000000; ec = 1; end
        16'b0001011000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001011000000000; ec = 1; end
        16'b0010110000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010110000000000; ec = 1; end
        16'b0101100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000101100000000000; ec = 1; end
        16'b1011000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001011000000000000; ec = 1; end
        16'b1110110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010110000000000000; ec = 1; end
        16'b0101011000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000101100000000000000; ec = 1; end
        16'b1010110001101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001011000000000000000; ec = 1; end
        16'b1101010100110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010110000000000000000; ec = 1; end
        16'b0010011110001111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000101100000000000000000; ec = 1; end
        16'b0100111100011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001011000000000000000000; ec = 1; end
        16'b1001111000111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010110000000000000000000; ec = 1; end
        16'b1011000110010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000101100000000000000000000; ec = 1; end
        16'b1110111011000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001011000000000000000000000; ec = 1; end
        16'b0101000001100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010110000000000000000000000; ec = 1; end
        16'b1010000011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000101100000000000000000000000; ec = 1; end
        16'b1100110001100001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001011000000000000000000000000; ec = 1; end
        16'b0001010100101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010110000000000000000000000000; ec = 1; end
        16'b0010101001011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000101100000000000000000000000000; ec = 1; end
        16'b0101010010111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001011000000000000000000000000000; ec = 1; end
        16'b1010100101111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010110000000000000000000000000000; ec = 1; end
        16'b1101111100011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000101100000000000000000000000000000; ec = 1; end
        16'b0011001111010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000001011000000000000000000000000000000; ec = 1; end
        16'b0110011110101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000010110000000000000000000000000000000; ec = 1; end
        16'b1100111101011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000101100000000000000000000000000000000; ec = 1; end
        16'b0001001101010101:begin data = code ^ 80'b00000000000000000000000000000000000000000001011000000000000000000000000000000000; ec = 1; end
        16'b0010011010101010:begin data = code ^ 80'b00000000000000000000000000000000000000000010110000000000000000000000000000000000; ec = 1; end
        16'b0100110101010100:begin data = code ^ 80'b00000000000000000000000000000000000000000101100000000000000000000000000000000000; ec = 1; end
        16'b1001101010101000:begin data = code ^ 80'b00000000000000000000000000000000000000001011000000000000000000000000000000000000; ec = 1; end
        16'b1011100010111101:begin data = code ^ 80'b00000000000000000000000000000000000000010110000000000000000000000000000000000000; ec = 1; end
        16'b1111110010010111:begin data = code ^ 80'b00000000000000000000000000000000000000101100000000000000000000000000000000000000; ec = 1; end
        16'b0111010011000011:begin data = code ^ 80'b00000000000000000000000000000000000001011000000000000000000000000000000000000000; ec = 1; end
        16'b1110100110000110:begin data = code ^ 80'b00000000000000000000000000000000000010110000000000000000000000000000000000000000; ec = 1; end
        16'b0101111011100001:begin data = code ^ 80'b00000000000000000000000000000000000101100000000000000000000000000000000000000000; ec = 1; end
        16'b1011110111000010:begin data = code ^ 80'b00000000000000000000000000000000001011000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011001101001:begin data = code ^ 80'b00000000000000000000000000000000010110000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000100111111:begin data = code ^ 80'b00000000000000000000000000000000101100000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001001111110:begin data = code ^ 80'b00000000000000000000000000000001011000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100100010001:begin data = code ^ 80'b00000000000000000000000000000010110000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001000100010:begin data = code ^ 80'b00000000000000000000000000000101100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010010001000100:begin data = code ^ 80'b00000000000000000000000000001011000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100010001000:begin data = code ^ 80'b00000000000000000000000000010110000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000100010000:begin data = code ^ 80'b00000000000000000000000000101100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111111001101:begin data = code ^ 80'b00000000000000000000000001011000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101001001110111:begin data = code ^ 80'b00000000000000000000000010110000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010100100000011:begin data = code ^ 80'b00000000000000000000000101100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101001000000110:begin data = code ^ 80'b00000000000000000000001011000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010010000001100:begin data = code ^ 80'b00000000000000000000010110000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100010111110101:begin data = code ^ 80'b00000000000000000000101100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011000000111:begin data = code ^ 80'b00000000000000000001011000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000110000001110:begin data = code ^ 80'b00000000000000000010110000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100000011100:begin data = code ^ 80'b00000000000000000101100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000000111000:begin data = code ^ 80'b00000000000000001011000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000001110000:begin data = code ^ 80'b00000000000000010110000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100000011100000:begin data = code ^ 80'b00000000000000101100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000110000101101:begin data = code ^ 80'b00000000000001011000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100001011010:begin data = code ^ 80'b00000000000010110000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000010110100:begin data = code ^ 80'b00000000000101100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000101101000:begin data = code ^ 80'b00000000001011000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001011010000:begin data = code ^ 80'b00000000010110000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100001001101:begin data = code ^ 80'b00000000101100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000010011010:begin data = code ^ 80'b00000001011000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000100110100:begin data = code ^ 80'b00000010110000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001001101000:begin data = code ^ 80'b00000101100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010011010000:begin data = code ^ 80'b00001011000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010001001101:begin data = code ^ 80'b00010110000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010101110111:begin data = code ^ 80'b00101100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011100000011:begin data = code ^ 80'b01011000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000001111101011:begin data = code ^ 80'b10110000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000000001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001101; ec = 1; end
        16'b0000000000011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000011010; ec = 1; end
        16'b0000000000110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110100; ec = 1; end
        16'b0000000001101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001101000; ec = 1; end
        16'b0000000011010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000011010000; ec = 1; end
        16'b0000000110100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000110100000; ec = 1; end
        16'b0000001101000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001101000000; ec = 1; end
        16'b0000011010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000011010000000; ec = 1; end
        16'b0000110100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000110100000000; ec = 1; end
        16'b0001101000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001101000000000; ec = 1; end
        16'b0011010000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000011010000000000; ec = 1; end
        16'b0110100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000110100000000000; ec = 1; end
        16'b1101000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001101000000000000; ec = 1; end
        16'b0010110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000011010000000000000; ec = 1; end
        16'b0101101111011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000110100000000000000; ec = 1; end
        16'b1011011110110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001101000000000000000; ec = 1; end
        16'b1110001010000101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000011010000000000000000; ec = 1; end
        16'b0100100011100111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000110100000000000000000; ec = 1; end
        16'b1001000111001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001101000000000000000000; ec = 1; end
        16'b1010111001110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000011010000000000000000000; ec = 1; end
        16'b1101000100001111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000110100000000000000000000; ec = 1; end
        16'b0010111111110011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001101000000000000000000000; ec = 1; end
        16'b0101111111100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000011010000000000000000000000; ec = 1; end
        16'b1011111111001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000110100000000000000000000000; ec = 1; end
        16'b1111001001110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001101000000000000000000000000; ec = 1; end
        16'b0110100100000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000011010000000000000000000000000; ec = 1; end
        16'b1101001000001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000110100000000000000000000000000; ec = 1; end
        16'b0010100111110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001101000000000000000000000000000; ec = 1; end
        16'b0101001111100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000011010000000000000000000000000000; ec = 1; end
        16'b1010011111000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000110100000000000000000000000000000; ec = 1; end
        16'b1100001001100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001101000000000000000000000000000000; ec = 1; end
        16'b0000100100100111:begin data = code ^ 80'b00000000000000000000000000000000000000000000011010000000000000000000000000000000; ec = 1; end
        16'b0001001001001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000110100000000000000000000000000000000; ec = 1; end
        16'b0010010010011100:begin data = code ^ 80'b00000000000000000000000000000000000000000001101000000000000000000000000000000000; ec = 1; end
        16'b0100100100111000:begin data = code ^ 80'b00000000000000000000000000000000000000000011010000000000000000000000000000000000; ec = 1; end
        16'b1001001001110000:begin data = code ^ 80'b00000000000000000000000000000000000000000110100000000000000000000000000000000000; ec = 1; end
        16'b1010100100001101:begin data = code ^ 80'b00000000000000000000000000000000000000001101000000000000000000000000000000000000; ec = 1; end
        16'b1101111111110111:begin data = code ^ 80'b00000000000000000000000000000000000000011010000000000000000000000000000000000000; ec = 1; end
        16'b0011001000000011:begin data = code ^ 80'b00000000000000000000000000000000000000110100000000000000000000000000000000000000; ec = 1; end
        16'b0110010000000110:begin data = code ^ 80'b00000000000000000000000000000000000001101000000000000000000000000000000000000000; ec = 1; end
        16'b1100100000001100:begin data = code ^ 80'b00000000000000000000000000000000000011010000000000000000000000000000000000000000; ec = 1; end
        16'b0001110111110101:begin data = code ^ 80'b00000000000000000000000000000000000110100000000000000000000000000000000000000000; ec = 1; end
        16'b0011101111101010:begin data = code ^ 80'b00000000000000000000000000000000001101000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011111010100:begin data = code ^ 80'b00000000000000000000000000000000011010000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111110101000:begin data = code ^ 80'b00000000000000000000000000000000110100000000000000000000000000000000000000000000; ec = 1; end
        16'b0101001010111101:begin data = code ^ 80'b00000000000000000000000000000001101000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010010101111010:begin data = code ^ 80'b00000000000000000000000000000011010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011100011001:begin data = code ^ 80'b00000000000000000000000000000110100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001111011111:begin data = code ^ 80'b00000000000000000000000000001101000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011110111110:begin data = code ^ 80'b00000000000000000000000000011010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111101111100:begin data = code ^ 80'b00000000000000000000000000110100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001111011111000:begin data = code ^ 80'b00000000000000000000000001101000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011110111110000:begin data = code ^ 80'b00000000000000000000000011010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111101111100000:begin data = code ^ 80'b00000000000000000000000110100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011111000000:begin data = code ^ 80'b00000000000000000000001101000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001001101101:begin data = code ^ 80'b00000000000000000000011010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100010011011010:begin data = code ^ 80'b00000000000000000000110100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000010001011001:begin data = code ^ 80'b00000000000000000001101000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100010110010:begin data = code ^ 80'b00000000000000000011010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000101100100:begin data = code ^ 80'b00000000000000000110100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010001011001000:begin data = code ^ 80'b00000000000000001101000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100010110010000:begin data = code ^ 80'b00000000000000011010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101100100000:begin data = code ^ 80'b00000000000000110100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001101110101101:begin data = code ^ 80'b00000000000001101000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011101010110111:begin data = code ^ 80'b00000000000011010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100010000011:begin data = code ^ 80'b00000000000110100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111110011101011:begin data = code ^ 80'b00000000001101000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100111010110:begin data = code ^ 80'b00000000011010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111001000001:begin data = code ^ 80'b00000000110100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111110010000010:begin data = code ^ 80'b00000001101000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111010011101001:begin data = code ^ 80'b00000011010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110100111010010:begin data = code ^ 80'b00000110100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111001001001:begin data = code ^ 80'b00001101000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110010010010:begin data = code ^ 80'b00011010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111010011001001:begin data = code ^ 80'b00110100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110010001111111:begin data = code ^ 80'b01101000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100011111110:begin data = code ^ 80'b11010000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000000001111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001111; ec = 1; end
        16'b0000000000011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000011110; ec = 1; end
        16'b0000000000111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000111100; ec = 1; end
        16'b0000000001111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001111000; ec = 1; end
        16'b0000000011110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000011110000; ec = 1; end
        16'b0000000111100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000111100000; ec = 1; end
        16'b0000001111000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001111000000; ec = 1; end
        16'b0000011110000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000011110000000; ec = 1; end
        16'b0000111100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000111100000000; ec = 1; end
        16'b0001111000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001111000000000; ec = 1; end
        16'b0011110000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000011110000000000; ec = 1; end
        16'b0111100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000111100000000000; ec = 1; end
        16'b1111000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001111000000000000; ec = 1; end
        16'b0110110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000011110000000000000; ec = 1; end
        16'b1101101111011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000111100000000000000; ec = 1; end
        16'b0011101001011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001111000000000000000; ec = 1; end
        16'b0111010010110010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000011110000000000000000; ec = 1; end
        16'b1110100101100100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000111100000000000000000; ec = 1; end
        16'b0101111100100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001111000000000000000000; ec = 1; end
        16'b1011111001001010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000011110000000000000000000; ec = 1; end
        16'b1111000101111001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000111100000000000000000000; ec = 1; end
        16'b0110111100011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001111000000000000000000000; ec = 1; end
        16'b1101111000111110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000011110000000000000000000000; ec = 1; end
        16'b0011000110010001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000111100000000000000000000000; ec = 1; end
        16'b0110001100100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001111000000000000000000000000; ec = 1; end
        16'b1100011001000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000011110000000000000000000000000; ec = 1; end
        16'b0000000101100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000111100000000000000000000000000; ec = 1; end
        16'b0000001011001010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001111000000000000000000000000000; ec = 1; end
        16'b0000010110010100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000011110000000000000000000000000000; ec = 1; end
        16'b0000101100101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000111100000000000000000000000000000; ec = 1; end
        16'b0001011001010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000001111000000000000000000000000000000; ec = 1; end
        16'b0010110010100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000011110000000000000000000000000000000; ec = 1; end
        16'b0101100101000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000111100000000000000000000000000000000; ec = 1; end
        16'b1011001010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000001111000000000000000000000000000000000; ec = 1; end
        16'b1110100011101101:begin data = code ^ 80'b00000000000000000000000000000000000000000011110000000000000000000000000000000000; ec = 1; end
        16'b0101110000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000111100000000000000000000000000000000000; ec = 1; end
        16'b1011100001101110:begin data = code ^ 80'b00000000000000000000000000000000000000001111000000000000000000000000000000000000; ec = 1; end
        16'b1111110100110001:begin data = code ^ 80'b00000000000000000000000000000000000000011110000000000000000000000000000000000000; ec = 1; end
        16'b0111011110001111:begin data = code ^ 80'b00000000000000000000000000000000000000111100000000000000000000000000000000000000; ec = 1; end
        16'b1110111100011110:begin data = code ^ 80'b00000000000000000000000000000000000001111000000000000000000000000000000000000000; ec = 1; end
        16'b0101001111010001:begin data = code ^ 80'b00000000000000000000000000000000000011110000000000000000000000000000000000000000; ec = 1; end
        16'b1010011110100010:begin data = code ^ 80'b00000000000000000000000000000000000111100000000000000000000000000000000000000000; ec = 1; end
        16'b1100001010101001:begin data = code ^ 80'b00000000000000000000000000000000001111000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100010111111:begin data = code ^ 80'b00000000000000000000000000000000011110000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000101111110:begin data = code ^ 80'b00000000000000000000000000000000111100000000000000000000000000000000000000000000; ec = 1; end
        16'b0010001011111100:begin data = code ^ 80'b00000000000000000000000000000001111000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100010111111000:begin data = code ^ 80'b00000000000000000000000000000011110000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101111110000:begin data = code ^ 80'b00000000000000000000000000000111100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001101000001101:begin data = code ^ 80'b00000000000000000000000000001111000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011100111110111:begin data = code ^ 80'b00000000000000000000000000011110000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111000000011:begin data = code ^ 80'b00000000000000000000000000111100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000111101011:begin data = code ^ 80'b00000000000000000000000001111000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001111010110:begin data = code ^ 80'b00000000000000000000000011110000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100101001000001:begin data = code ^ 80'b00000000000000000000000111100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001010010000010:begin data = code ^ 80'b00000000000000000000001111000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010010011101001:begin data = code ^ 80'b00000000000000000000011110000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100010000111111:begin data = code ^ 80'b00000000000000000000111100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000010110010011:begin data = code ^ 80'b00000000000000000001111000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101100100110:begin data = code ^ 80'b00000000000000000011110000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011001001100:begin data = code ^ 80'b00000000000000000111100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110010011000:begin data = code ^ 80'b00000000000000001111000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101100100110000:begin data = code ^ 80'b00000000000000011110000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011001001100000:begin data = code ^ 80'b00000000000000111100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110100100101101:begin data = code ^ 80'b00000000000001111000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111110110111:begin data = code ^ 80'b00000000000011110000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111101101110:begin data = code ^ 80'b00000000000111100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111001100110001:begin data = code ^ 80'b00000000001111000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110101110001111:begin data = code ^ 80'b00000000011110000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101011100011110:begin data = code ^ 80'b00000000111100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010001111010001:begin data = code ^ 80'b00000001111000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011110100010:begin data = code ^ 80'b00000011110000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111101000100:begin data = code ^ 80'b00000111100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001101100101:begin data = code ^ 80'b00001111000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010101100100111:begin data = code ^ 80'b00011110000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101101110100011:begin data = code ^ 80'b00111100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011101010101011:begin data = code ^ 80'b01111000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111010101010110:begin data = code ^ 80'b11110000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000000000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000011; ec = 1; end
        16'b0000000000000101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000101; ec = 1; end
        16'b0000000000000110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000110; ec = 1; end
        16'b0000000000001001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001001; ec = 1; end
        16'b0000000000001010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001010; ec = 1; end
        16'b0000000000001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000001100; ec = 1; end
        16'b0000000000010001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010001; ec = 1; end
        16'b0000000000010010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010010; ec = 1; end
        16'b0000000000010100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000010100; ec = 1; end
        16'b0000000000011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000011000; ec = 1; end
        16'b0000000000100001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100001; ec = 1; end
        16'b0000000000100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100010; ec = 1; end
        16'b0000000000100100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000100100; ec = 1; end
        16'b0000000000101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000101000; ec = 1; end
        16'b0000000000110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000000110000; ec = 1; end
        16'b0000000001000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000001; ec = 1; end
        16'b0000000001000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000010; ec = 1; end
        16'b0000000001000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001000100; ec = 1; end
        16'b0000000001001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001001000; ec = 1; end
        16'b0000000001010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001010000; ec = 1; end
        16'b0000000001100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000001100000; ec = 1; end
        16'b0000000010000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000001; ec = 1; end
        16'b0000000010000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000010; ec = 1; end
        16'b0000000010000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010000100; ec = 1; end
        16'b0000000010001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010001000; ec = 1; end
        16'b0000000010010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010010000; ec = 1; end
        16'b0000000010100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000010100000; ec = 1; end
        16'b0000000011000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000011000000; ec = 1; end
        16'b0000000100000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100000001; ec = 1; end
        16'b0000000100000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100000010; ec = 1; end
        16'b0000000100000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100000100; ec = 1; end
        16'b0000000100001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100001000; ec = 1; end
        16'b0000000100010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100010000; ec = 1; end
        16'b0000000100100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000100100000; ec = 1; end
        16'b0000000101000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000101000000; ec = 1; end
        16'b0000000110000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000000110000000; ec = 1; end
        16'b0000001000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000000001; ec = 1; end
        16'b0000001000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000000010; ec = 1; end
        16'b0000001000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000000100; ec = 1; end
        16'b0000001000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000001000; ec = 1; end
        16'b0000001000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000010000; ec = 1; end
        16'b0000001000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001000100000; ec = 1; end
        16'b0000001001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001001000000; ec = 1; end
        16'b0000001010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001010000000; ec = 1; end
        16'b0000001100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000001100000000; ec = 1; end
        16'b0000010000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000000001; ec = 1; end
        16'b0000010000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000000010; ec = 1; end
        16'b0000010000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000000100; ec = 1; end
        16'b0000010000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000001000; ec = 1; end
        16'b0000010000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000010000; ec = 1; end
        16'b0000010000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010000100000; ec = 1; end
        16'b0000010001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010001000000; ec = 1; end
        16'b0000010010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010010000000; ec = 1; end
        16'b0000010100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000010100000000; ec = 1; end
        16'b0000011000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000011000000000; ec = 1; end
        16'b0000100000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000001; ec = 1; end
        16'b0000100000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000010; ec = 1; end
        16'b0000100000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000000100; ec = 1; end
        16'b0000100000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000001000; ec = 1; end
        16'b0000100000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000010000; ec = 1; end
        16'b0000100000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100000100000; ec = 1; end
        16'b0000100001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100001000000; ec = 1; end
        16'b0000100010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100010000000; ec = 1; end
        16'b0000100100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000100100000000; ec = 1; end
        16'b0000101000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000101000000000; ec = 1; end
        16'b0000110000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000000110000000000; ec = 1; end
        16'b0001000000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000001; ec = 1; end
        16'b0001000000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000010; ec = 1; end
        16'b0001000000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000000100; ec = 1; end
        16'b0001000000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000001000; ec = 1; end
        16'b0001000000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000010000; ec = 1; end
        16'b0001000000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000000100000; ec = 1; end
        16'b0001000001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000001000000; ec = 1; end
        16'b0001000010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000010000000; ec = 1; end
        16'b0001000100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001000100000000; ec = 1; end
        16'b0001001000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001001000000000; ec = 1; end
        16'b0001010000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001010000000000; ec = 1; end
        16'b0001100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000001100000000000; ec = 1; end
        16'b0010000000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000001; ec = 1; end
        16'b0010000000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000010; ec = 1; end
        16'b0010000000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000000100; ec = 1; end
        16'b0010000000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000001000; ec = 1; end
        16'b0010000000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000010000; ec = 1; end
        16'b0010000000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000000100000; ec = 1; end
        16'b0010000001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000001000000; ec = 1; end
        16'b0010000010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000010000000; ec = 1; end
        16'b0010000100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010000100000000; ec = 1; end
        16'b0010001000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010001000000000; ec = 1; end
        16'b0010010000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010010000000000; ec = 1; end
        16'b0010100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000010100000000000; ec = 1; end
        16'b0011000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000011000000000000; ec = 1; end
        16'b0100000000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000001; ec = 1; end
        16'b0100000000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000010; ec = 1; end
        16'b0100000000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000000100; ec = 1; end
        16'b0100000000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000001000; ec = 1; end
        16'b0100000000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000010000; ec = 1; end
        16'b0100000000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000000100000; ec = 1; end
        16'b0100000001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000001000000; ec = 1; end
        16'b0100000010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000010000000; ec = 1; end
        16'b0100000100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100000100000000; ec = 1; end
        16'b0100001000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100001000000000; ec = 1; end
        16'b0100010000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100010000000000; ec = 1; end
        16'b0100100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000100100000000000; ec = 1; end
        16'b0101000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000101000000000000; ec = 1; end
        16'b0110000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000000110000000000000; ec = 1; end
        16'b1000000000000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000001; ec = 1; end
        16'b1000000000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000010; ec = 1; end
        16'b1000000000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000000100; ec = 1; end
        16'b1000000000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000001000; ec = 1; end
        16'b1000000000010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000010000; ec = 1; end
        16'b1000000000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000000100000; ec = 1; end
        16'b1000000001000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000001000000; ec = 1; end
        16'b1000000010000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000010000000; ec = 1; end
        16'b1000000100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000000100000000; ec = 1; end
        16'b1000001000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000001000000000; ec = 1; end
        16'b1000010000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000010000000000; ec = 1; end
        16'b1000100000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001000100000000000; ec = 1; end
        16'b1001000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001001000000000000; ec = 1; end
        16'b1010000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001010000000000000; ec = 1; end
        16'b1100000000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000001100000000000000; ec = 1; end
        16'b1000110111101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000001; ec = 1; end
        16'b1000110111101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000010; ec = 1; end
        16'b1000110111101001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000000100; ec = 1; end
        16'b1000110111100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000001000; ec = 1; end
        16'b1000110111111101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000010000; ec = 1; end
        16'b1000110111001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000000100000; ec = 1; end
        16'b1000110110101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000001000000; ec = 1; end
        16'b1000110101101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000010000000; ec = 1; end
        16'b1000110011101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000000100000000; ec = 1; end
        16'b1000111111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000001000000000; ec = 1; end
        16'b1000100111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000010000000000; ec = 1; end
        16'b1000010111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010000100000000000; ec = 1; end
        16'b1001110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010001000000000000; ec = 1; end
        16'b1010110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010010000000000000; ec = 1; end
        16'b1100110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000010100000000000000; ec = 1; end
        16'b0000110111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000011000000000000000; ec = 1; end
        16'b1001011000110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000000001; ec = 1; end
        16'b1001011000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000000010; ec = 1; end
        16'b1001011000110011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000000100; ec = 1; end
        16'b1001011000111111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000001000; ec = 1; end
        16'b1001011000100111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000010000; ec = 1; end
        16'b1001011000010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000000100000; ec = 1; end
        16'b1001011001110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000001000000; ec = 1; end
        16'b1001011010110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000010000000; ec = 1; end
        16'b1001011100110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000000100000000; ec = 1; end
        16'b1001010000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000001000000000; ec = 1; end
        16'b1001001000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000010000000000; ec = 1; end
        16'b1001111000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100000100000000000; ec = 1; end
        16'b1000011000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100001000000000000; ec = 1; end
        16'b1011011000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100010000000000000; ec = 1; end
        16'b1101011000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000100100000000000000; ec = 1; end
        16'b0001011000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000101000000000000000; ec = 1; end
        16'b0001101111011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000000110000000000000000; ec = 1; end
        16'b1010000110000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000000001; ec = 1; end
        16'b1010000110000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000000010; ec = 1; end
        16'b1010000110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000000100; ec = 1; end
        16'b1010000110001011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000001000; ec = 1; end
        16'b1010000110010011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000010000; ec = 1; end
        16'b1010000110100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000000100000; ec = 1; end
        16'b1010000111000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000001000000; ec = 1; end
        16'b1010000100000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000010000000; ec = 1; end
        16'b1010000010000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000000100000000; ec = 1; end
        16'b1010001110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000001000000000; ec = 1; end
        16'b1010010110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000010000000000; ec = 1; end
        16'b1010100110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000000100000000000; ec = 1; end
        16'b1011000110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000001000000000000; ec = 1; end
        16'b1000000110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000010000000000000; ec = 1; end
        16'b1110000110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001000100000000000000; ec = 1; end
        16'b0010000110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001001000000000000000; ec = 1; end
        16'b0010110001101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001010000000000000000; ec = 1; end
        16'b0011011110110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000001100000000000000000; ec = 1; end
        16'b1100111011101010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000000001; ec = 1; end
        16'b1100111011101001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000000010; ec = 1; end
        16'b1100111011101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000000100; ec = 1; end
        16'b1100111011100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000001000; ec = 1; end
        16'b1100111011111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000010000; ec = 1; end
        16'b1100111011001011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000000100000; ec = 1; end
        16'b1100111010101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000001000000; ec = 1; end
        16'b1100111001101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000010000000; ec = 1; end
        16'b1100111111101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000000100000000; ec = 1; end
        16'b1100110011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000001000000000; ec = 1; end
        16'b1100101011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000010000000000; ec = 1; end
        16'b1100011011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000000100000000000; ec = 1; end
        16'b1101111011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000001000000000000; ec = 1; end
        16'b1110111011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000010000000000000; ec = 1; end
        16'b1000111011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010000100000000000000; ec = 1; end
        16'b0100111011101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010001000000000000000; ec = 1; end
        16'b0100001100000110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010010000000000000000; ec = 1; end
        16'b0101100011011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000010100000000000000000; ec = 1; end
        16'b0110111101101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000011000000000000000000; ec = 1; end
        16'b0001000000111010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000000001; ec = 1; end
        16'b0001000000111001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000000010; ec = 1; end
        16'b0001000000111111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000000100; ec = 1; end
        16'b0001000000110011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000001000; ec = 1; end
        16'b0001000000101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000010000; ec = 1; end
        16'b0001000000011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000000100000; ec = 1; end
        16'b0001000001111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000001000000; ec = 1; end
        16'b0001000010111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000010000000; ec = 1; end
        16'b0001000100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000000100000000; ec = 1; end
        16'b0001001000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000001000000000; ec = 1; end
        16'b0001010000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000010000000000; ec = 1; end
        16'b0001100000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000000100000000000; ec = 1; end
        16'b0000000000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000001000000000000; ec = 1; end
        16'b0011000000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000010000000000000; ec = 1; end
        16'b0101000000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100000100000000000000; ec = 1; end
        16'b1001000000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100001000000000000000; ec = 1; end
        16'b1001110111010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100010000000000000000; ec = 1; end
        16'b1000011000001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000100100000000000000000; ec = 1; end
        16'b1011000110111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000101000000000000000000; ec = 1; end
        16'b1101111011010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000000110000000000000000000; ec = 1; end
        16'b0010000001110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000000001; ec = 1; end
        16'b0010000001110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000000010; ec = 1; end
        16'b0010000001110010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000000100; ec = 1; end
        16'b0010000001111110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000001000; ec = 1; end
        16'b0010000001100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000010000; ec = 1; end
        16'b0010000001010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000000100000; ec = 1; end
        16'b0010000000110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000001000000; ec = 1; end
        16'b0010000011110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000010000000; ec = 1; end
        16'b0010000101110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000000100000000; ec = 1; end
        16'b0010001001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000001000000000; ec = 1; end
        16'b0010010001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000010000000000; ec = 1; end
        16'b0010100001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000000100000000000; ec = 1; end
        16'b0011000001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000001000000000000; ec = 1; end
        16'b0000000001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000010000000000000; ec = 1; end
        16'b0110000001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000000100000000000000; ec = 1; end
        16'b1010000001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000001000000000000000; ec = 1; end
        16'b1010110110011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000010000000000000000; ec = 1; end
        16'b1011011001000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001000100000000000000000; ec = 1; end
        16'b1000000111110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001001000000000000000000; ec = 1; end
        16'b1110111010011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001010000000000000000000; ec = 1; end
        16'b0011000001001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000001100000000000000000000; ec = 1; end
        16'b0100000011101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000000001; ec = 1; end
        16'b0100000011101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000000010; ec = 1; end
        16'b0100000011101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000000100; ec = 1; end
        16'b0100000011100100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000001000; ec = 1; end
        16'b0100000011111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000010000; ec = 1; end
        16'b0100000011001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000000100000; ec = 1; end
        16'b0100000010101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000001000000; ec = 1; end
        16'b0100000001101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000010000000; ec = 1; end
        16'b0100000111101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000000100000000; ec = 1; end
        16'b0100001011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000001000000000; ec = 1; end
        16'b0100010011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000010000000000; ec = 1; end
        16'b0100100011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000000100000000000; ec = 1; end
        16'b0101000011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000001000000000000; ec = 1; end
        16'b0110000011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000010000000000000; ec = 1; end
        16'b0000000011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000000100000000000000; ec = 1; end
        16'b1100000011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000001000000000000000; ec = 1; end
        16'b1100110100000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000010000000000000000; ec = 1; end
        16'b1101011011011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010000100000000000000000; ec = 1; end
        16'b1110000101101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010001000000000000000000; ec = 1; end
        16'b1000111000000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010010000000000000000000; ec = 1; end
        16'b0101000011010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000010100000000000000000000; ec = 1; end
        16'b0110000010011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000011000000000000000000000; ec = 1; end
        16'b1000000111011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000000001; ec = 1; end
        16'b1000000111011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000000010; ec = 1; end
        16'b1000000111011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000000100; ec = 1; end
        16'b1000000111010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000001000; ec = 1; end
        16'b1000000111001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000010000; ec = 1; end
        16'b1000000111111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000000100000; ec = 1; end
        16'b1000000110011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000001000000; ec = 1; end
        16'b1000000101011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000010000000; ec = 1; end
        16'b1000000011011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000000100000000; ec = 1; end
        16'b1000001111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000001000000000; ec = 1; end
        16'b1000010111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000010000000000; ec = 1; end
        16'b1000100111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000000100000000000; ec = 1; end
        16'b1001000111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000001000000000000; ec = 1; end
        16'b1010000111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000010000000000000; ec = 1; end
        16'b1100000111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000000100000000000000; ec = 1; end
        16'b0000000111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000001000000000000000; ec = 1; end
        16'b0000110000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000010000000000000000; ec = 1; end
        16'b0001011111101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100000100000000000000000; ec = 1; end
        16'b0010000001011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100001000000000000000000; ec = 1; end
        16'b0100111100110011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100010000000000000000000; ec = 1; end
        16'b1001000111100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000100100000000000000000000; ec = 1; end
        16'b1010000110101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000101000000000000000000000; ec = 1; end
        16'b1100000100110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000000110000000000000000000000; ec = 1; end
        16'b1000111001011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000000001; ec = 1; end
        16'b1000111001011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000000010; ec = 1; end
        16'b1000111001011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000000100; ec = 1; end
        16'b1000111001010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000001000; ec = 1; end
        16'b1000111001001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000010000; ec = 1; end
        16'b1000111001111101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000000100000; ec = 1; end
        16'b1000111000011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000001000000; ec = 1; end
        16'b1000111011011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000010000000; ec = 1; end
        16'b1000111101011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000000100000000; ec = 1; end
        16'b1000110001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000001000000000; ec = 1; end
        16'b1000101001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000010000000000; ec = 1; end
        16'b1000011001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000000100000000000; ec = 1; end
        16'b1001111001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000001000000000000; ec = 1; end
        16'b1010111001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000010000000000000; ec = 1; end
        16'b1100111001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000000100000000000000; ec = 1; end
        16'b0000111001011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000001000000000000000; ec = 1; end
        16'b0000001110110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000010000000000000000; ec = 1; end
        16'b0001100001101010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000000100000000000000000; ec = 1; end
        16'b0010111111011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000001000000000000000000; ec = 1; end
        16'b0100000010110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000010000000000000000000; ec = 1; end
        16'b1001111001100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001000100000000000000000000; ec = 1; end
        16'b1010111000101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001001000000000000000000000; ec = 1; end
        16'b1100111010110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001010000000000000000000000; ec = 1; end
        16'b0000111110000101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000001100000000000000000000000; ec = 1; end
        16'b1001000101010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000000001; ec = 1; end
        16'b1001000101010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000000010; ec = 1; end
        16'b1001000101010011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000000100; ec = 1; end
        16'b1001000101011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000001000; ec = 1; end
        16'b1001000101000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000010000; ec = 1; end
        16'b1001000101110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000000100000; ec = 1; end
        16'b1001000100010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000001000000; ec = 1; end
        16'b1001000111010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000010000000; ec = 1; end
        16'b1001000001010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000000100000000; ec = 1; end
        16'b1001001101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000001000000000; ec = 1; end
        16'b1001010101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000010000000000; ec = 1; end
        16'b1001100101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000000100000000000; ec = 1; end
        16'b1000000101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000001000000000000; ec = 1; end
        16'b1011000101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000010000000000000; ec = 1; end
        16'b1101000101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000000100000000000000; ec = 1; end
        16'b0001000101010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000001000000000000000; ec = 1; end
        16'b0001110010111010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000010000000000000000; ec = 1; end
        16'b0000011101100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000000100000000000000000; ec = 1; end
        16'b0011000011010100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000001000000000000000000; ec = 1; end
        16'b0101111110111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000010000000000000000000; ec = 1; end
        16'b1000000101101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010000100000000000000000000; ec = 1; end
        16'b1011000100100001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010001000000000000000000000; ec = 1; end
        16'b1101000110111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010010000000000000000000000; ec = 1; end
        16'b0001000010001111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000010100000000000000000000000; ec = 1; end
        16'b0001111100001010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000011000000000000000000000000; ec = 1; end
        16'b1010111101000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000000001; ec = 1; end
        16'b1010111101000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000000010; ec = 1; end
        16'b1010111101000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000000100; ec = 1; end
        16'b1010111101001011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000001000; ec = 1; end
        16'b1010111101010011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000010000; ec = 1; end
        16'b1010111101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000000100000; ec = 1; end
        16'b1010111100000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000001000000; ec = 1; end
        16'b1010111111000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000010000000; ec = 1; end
        16'b1010111001000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000000100000000; ec = 1; end
        16'b1010110101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000001000000000; ec = 1; end
        16'b1010101101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000010000000000; ec = 1; end
        16'b1010011101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000000100000000000; ec = 1; end
        16'b1011111101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000001000000000000; ec = 1; end
        16'b1000111101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000010000000000000; ec = 1; end
        16'b1110111101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000000100000000000000; ec = 1; end
        16'b0010111101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000001000000000000000; ec = 1; end
        16'b0010001010101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000010000000000000000; ec = 1; end
        16'b0011100101110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000000100000000000000000; ec = 1; end
        16'b0000111011000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000001000000000000000000; ec = 1; end
        16'b0110000110101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000010000000000000000000; ec = 1; end
        16'b1011111101111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100000100000000000000000000; ec = 1; end
        16'b1000111100110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100001000000000000000000000; ec = 1; end
        16'b1110111110101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100010000000000000000000000; ec = 1; end
        16'b0010111010011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000100100000000000000000000000; ec = 1; end
        16'b0010000100011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000101000000000000000000000000; ec = 1; end
        16'b0011111000010100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000000110000000000000000000000000; ec = 1; end
        16'b1101001101101010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000000001; ec = 1; end
        16'b1101001101101001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000000010; ec = 1; end
        16'b1101001101101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000000100; ec = 1; end
        16'b1101001101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000001000; ec = 1; end
        16'b1101001101111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000010000; ec = 1; end
        16'b1101001101001011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000000100000; ec = 1; end
        16'b1101001100101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000001000000; ec = 1; end
        16'b1101001111101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000010000000; ec = 1; end
        16'b1101001001101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000000100000000; ec = 1; end
        16'b1101000101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000001000000000; ec = 1; end
        16'b1101011101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000010000000000; ec = 1; end
        16'b1101101101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000000100000000000; ec = 1; end
        16'b1100001101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000001000000000000; ec = 1; end
        16'b1111001101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000010000000000000; ec = 1; end
        16'b1001001101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000000100000000000000; ec = 1; end
        16'b0101001101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000001000000000000000; ec = 1; end
        16'b0101111010000110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000010000000000000000; ec = 1; end
        16'b0100010101011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000000100000000000000000; ec = 1; end
        16'b0111001011101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000001000000000000000000; ec = 1; end
        16'b0001110110000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000010000000000000000000; ec = 1; end
        16'b1100001101010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000000100000000000000000000; ec = 1; end
        16'b1111001100011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000001000000000000000000000; ec = 1; end
        16'b1001001110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000010000000000000000000000; ec = 1; end
        16'b0101001010110011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001000100000000000000000000000; ec = 1; end
        16'b0101110100110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001001000000000000000000000000; ec = 1; end
        16'b0100001000111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001010000000000000000000000000; ec = 1; end
        16'b0111110000101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000001100000000000000000000000000; ec = 1; end
        16'b0010101100111010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000000001; ec = 1; end
        16'b0010101100111001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000000010; ec = 1; end
        16'b0010101100111111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000000100; ec = 1; end
        16'b0010101100110011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000001000; ec = 1; end
        16'b0010101100101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000010000; ec = 1; end
        16'b0010101100011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000000100000; ec = 1; end
        16'b0010101101111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000001000000; ec = 1; end
        16'b0010101110111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000010000000; ec = 1; end
        16'b0010101000111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000000100000000; ec = 1; end
        16'b0010100100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000001000000000; ec = 1; end
        16'b0010111100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000010000000000; ec = 1; end
        16'b0010001100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000000100000000000; ec = 1; end
        16'b0011101100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000001000000000000; ec = 1; end
        16'b0000101100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000010000000000000; ec = 1; end
        16'b0110101100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000000100000000000000; ec = 1; end
        16'b1010101100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000001000000000000000; ec = 1; end
        16'b1010011011010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000010000000000000000; ec = 1; end
        16'b1011110100001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000000100000000000000000; ec = 1; end
        16'b1000101010111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000001000000000000000000; ec = 1; end
        16'b1110010111010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000010000000000000000000; ec = 1; end
        16'b0011101100000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000000100000000000000000000; ec = 1; end
        16'b0000101101001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000001000000000000000000000; ec = 1; end
        16'b0110101111010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000010000000000000000000000; ec = 1; end
        16'b1010101011100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010000100000000000000000000000; ec = 1; end
        16'b1010010101100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010001000000000000000000000000; ec = 1; end
        16'b1011101001101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010010000000000000000000000000; ec = 1; end
        16'b1000010001111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000010100000000000000000000000000; ec = 1; end
        16'b1111100001010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000011000000000000000000000000000; ec = 1; end
        16'b0101011001110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000000001; ec = 1; end
        16'b0101011001110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000000010; ec = 1; end
        16'b0101011001110010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000000100; ec = 1; end
        16'b0101011001111110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000001000; ec = 1; end
        16'b0101011001100110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000010000; ec = 1; end
        16'b0101011001010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000000100000; ec = 1; end
        16'b0101011000110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000001000000; ec = 1; end
        16'b0101011011110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000010000000; ec = 1; end
        16'b0101011101110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000000100000000; ec = 1; end
        16'b0101010001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000001000000000; ec = 1; end
        16'b0101001001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000010000000000; ec = 1; end
        16'b0101111001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000000100000000000; ec = 1; end
        16'b0100011001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000001000000000000; ec = 1; end
        16'b0111011001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000010000000000000; ec = 1; end
        16'b0001011001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000000100000000000000; ec = 1; end
        16'b1101011001110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000001000000000000000; ec = 1; end
        16'b1101101110011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000010000000000000000; ec = 1; end
        16'b1100000001000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000000100000000000000000; ec = 1; end
        16'b1111011111110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000001000000000000000000; ec = 1; end
        16'b1001100010011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000010000000000000000000; ec = 1; end
        16'b0100011001001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000000100000000000000000000; ec = 1; end
        16'b0111011000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000001000000000000000000000; ec = 1; end
        16'b0001011010011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000010000000000000000000000; ec = 1; end
        16'b1101011110101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100000100000000000000000000000; ec = 1; end
        16'b1101100000101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100001000000000000000000000000; ec = 1; end
        16'b1100011100100001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100010000000000000000000000000; ec = 1; end
        16'b1111100100110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000100100000000000000000000000000; ec = 1; end
        16'b1000010100011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000101000000000000000000000000000; ec = 1; end
        16'b0111110101001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000000110000000000000000000000000000; ec = 1; end
        16'b1010110011101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000000001; ec = 1; end
        16'b1010110011101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000000010; ec = 1; end
        16'b1010110011101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000000100; ec = 1; end
        16'b1010110011100100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000001000; ec = 1; end
        16'b1010110011111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000010000; ec = 1; end
        16'b1010110011001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000000100000; ec = 1; end
        16'b1010110010101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000001000000; ec = 1; end
        16'b1010110001101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000010000000; ec = 1; end
        16'b1010110111101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000000100000000; ec = 1; end
        16'b1010111011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000001000000000; ec = 1; end
        16'b1010100011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000010000000000; ec = 1; end
        16'b1010010011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000000100000000000; ec = 1; end
        16'b1011110011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000001000000000000; ec = 1; end
        16'b1000110011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000010000000000000; ec = 1; end
        16'b1110110011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000000100000000000000; ec = 1; end
        16'b0010110011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000001000000000000000; ec = 1; end
        16'b0010000100000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000010000000000000000; ec = 1; end
        16'b0011101011011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000000100000000000000000; ec = 1; end
        16'b0000110101101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000001000000000000000000; ec = 1; end
        16'b0110001000000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000010000000000000000000; ec = 1; end
        16'b1011110011010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000000100000000000000000000; ec = 1; end
        16'b1000110010011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000001000000000000000000000; ec = 1; end
        16'b1110110000000000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000010000000000000000000000; ec = 1; end
        16'b0010110100110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000000100000000000000000000000; ec = 1; end
        16'b0010001010110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000001000000000000000000000000; ec = 1; end
        16'b0011110110111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000010000000000000000000000000; ec = 1; end
        16'b0000001110101111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001000100000000000000000000000000; ec = 1; end
        16'b0111111110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001001000000000000000000000000000; ec = 1; end
        16'b1000011111010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001010000000000000000000000000000; ec = 1; end
        16'b1111101010011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000001100000000000000000000000000000; ec = 1; end
        16'b1101010000110100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000000001; ec = 1; end
        16'b1101010000110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000000010; ec = 1; end
        16'b1101010000110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000000100; ec = 1; end
        16'b1101010000111101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000001000; ec = 1; end
        16'b1101010000100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000010000; ec = 1; end
        16'b1101010000010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000000100000; ec = 1; end
        16'b1101010001110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000001000000; ec = 1; end
        16'b1101010010110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000010000000; ec = 1; end
        16'b1101010100110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000000100000000; ec = 1; end
        16'b1101011000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000001000000000; ec = 1; end
        16'b1101000000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000010000000000; ec = 1; end
        16'b1101110000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000000100000000000; ec = 1; end
        16'b1100010000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000001000000000000; ec = 1; end
        16'b1111010000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000010000000000000; ec = 1; end
        16'b1001010000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000000100000000000000; ec = 1; end
        16'b0101010000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000001000000000000000; ec = 1; end
        16'b0101100111011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000010000000000000000; ec = 1; end
        16'b0100001000000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000000100000000000000000; ec = 1; end
        16'b0111010110110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000001000000000000000000; ec = 1; end
        16'b0001101011011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000010000000000000000000; ec = 1; end
        16'b1100010000001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000000100000000000000000000; ec = 1; end
        16'b1111010001000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000001000000000000000000000; ec = 1; end
        16'b1001010011011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000010000000000000000000000; ec = 1; end
        16'b0101010111101101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000000100000000000000000000000; ec = 1; end
        16'b0101101001101000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000001000000000000000000000000; ec = 1; end
        16'b0100010101100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000010000000000000000000000000; ec = 1; end
        16'b0111101101110110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010000100000000000000000000000000; ec = 1; end
        16'b0000011101011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010001000000000000000000000000000; ec = 1; end
        16'b1111111100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010010000000000000000000000000000; ec = 1; end
        16'b1000001001000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000010100000000000000000000000000000; ec = 1; end
        16'b0111100011011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000011000000000000000000000000000000; ec = 1; end
        16'b0010010110000110:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000000001; ec = 1; end
        16'b0010010110000101:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000000010; ec = 1; end
        16'b0010010110000011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000000100; ec = 1; end
        16'b0010010110001111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000001000; ec = 1; end
        16'b0010010110010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000010000; ec = 1; end
        16'b0010010110100111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000000100000; ec = 1; end
        16'b0010010111000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000001000000; ec = 1; end
        16'b0010010100000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000010000000; ec = 1; end
        16'b0010010010000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000000100000000; ec = 1; end
        16'b0010011110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000001000000000; ec = 1; end
        16'b0010000110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000010000000000; ec = 1; end
        16'b0010110110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000000100000000000; ec = 1; end
        16'b0011010110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000001000000000000; ec = 1; end
        16'b0000010110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000010000000000000; ec = 1; end
        16'b0110010110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000000100000000000000; ec = 1; end
        16'b1010010110000111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000001000000000000000; ec = 1; end
        16'b1010100001101010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000010000000000000000; ec = 1; end
        16'b1011001110110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000000100000000000000000; ec = 1; end
        16'b1000010000000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000001000000000000000000; ec = 1; end
        16'b1110101101101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000010000000000000000000; ec = 1; end
        16'b0011010110111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000000100000000000000000000; ec = 1; end
        16'b0000010111110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000001000000000000000000000; ec = 1; end
        16'b0110010101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000010000000000000000000000; ec = 1; end
        16'b1010010001011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000000100000000000000000000000; ec = 1; end
        16'b1010101111011010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000001000000000000000000000000; ec = 1; end
        16'b1011010011010000:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000010000000000000000000000000; ec = 1; end
        16'b1000101011000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100000100000000000000000000000000; ec = 1; end
        16'b1111011011101100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100001000000000000000000000000000; ec = 1; end
        16'b0000111010111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100010000000000000000000000000000; ec = 1; end
        16'b0111001111110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000000100100000000000000000000000000000; ec = 1; end
        16'b1000100101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000000101000000000000000000000000000000; ec = 1; end
        16'b1111000110110010:begin data = code ^ 80'b00000000000000000000000000000000000000000000000110000000000000000000000000000000; ec = 1; end
        16'b0100101100001111:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000000001; ec = 1; end
        16'b0100101100001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000000010; ec = 1; end
        16'b0100101100001010:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000000100; ec = 1; end
        16'b0100101100000110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000001000; ec = 1; end
        16'b0100101100011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000010000; ec = 1; end
        16'b0100101100101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000000100000; ec = 1; end
        16'b0100101101001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000001000000; ec = 1; end
        16'b0100101110001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000010000000; ec = 1; end
        16'b0100101000001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000000100000000; ec = 1; end
        16'b0100100100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000001000000000; ec = 1; end
        16'b0100111100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000010000000000; ec = 1; end
        16'b0100001100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000000100000000000; ec = 1; end
        16'b0101101100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000001000000000000; ec = 1; end
        16'b0110101100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000010000000000000; ec = 1; end
        16'b0000101100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000000100000000000000; ec = 1; end
        16'b1100101100001110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000001000000000000000; ec = 1; end
        16'b1100011011100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000010000000000000000; ec = 1; end
        16'b1101110100111001:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000000100000000000000000; ec = 1; end
        16'b1110101010001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000001000000000000000000; ec = 1; end
        16'b1000010111100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000010000000000000000000; ec = 1; end
        16'b0101101100110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000000100000000000000000000; ec = 1; end
        16'b0110101101111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000001000000000000000000000; ec = 1; end
        16'b0000101111100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000010000000000000000000000; ec = 1; end
        16'b1100101011010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000000100000000000000000000000; ec = 1; end
        16'b1100010101010011:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000001000000000000000000000000; ec = 1; end
        16'b1101101001011001:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000010000000000000000000000000; ec = 1; end
        16'b1110010001001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000000100000000000000000000000000; ec = 1; end
        16'b1001100001100101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000001000000000000000000000000000; ec = 1; end
        16'b0110000000110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000010000000000000000000000000000; ec = 1; end
        16'b0001110101111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000001000100000000000000000000000000000; ec = 1; end
        16'b1110011111100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000001001000000000000000000000000000000; ec = 1; end
        16'b1001111100111011:begin data = code ^ 80'b00000000000000000000000000000000000000000000001010000000000000000000000000000000; ec = 1; end
        16'b0110111010001001:begin data = code ^ 80'b00000000000000000000000000000000000000000000001100000000000000000000000000000000; ec = 1; end
        16'b1001011000011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000000001; ec = 1; end
        16'b1001011000011110:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000000010; ec = 1; end
        16'b1001011000011000:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000000100; ec = 1; end
        16'b1001011000010100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000001000; ec = 1; end
        16'b1001011000001100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000010000; ec = 1; end
        16'b1001011000111100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000000100000; ec = 1; end
        16'b1001011001011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000001000000; ec = 1; end
        16'b1001011010011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000010000000; ec = 1; end
        16'b1001011100011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000000100000000; ec = 1; end
        16'b1001010000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000001000000000; ec = 1; end
        16'b1001001000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000010000000000; ec = 1; end
        16'b1001111000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000000100000000000; ec = 1; end
        16'b1000011000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000001000000000000; ec = 1; end
        16'b1011011000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000010000000000000; ec = 1; end
        16'b1101011000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000000100000000000000; ec = 1; end
        16'b0001011000011100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000001000000000000000; ec = 1; end
        16'b0001101111110001:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000010000000000000000; ec = 1; end
        16'b0000000000101011:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000000100000000000000000; ec = 1; end
        16'b0011011110011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000001000000000000000000; ec = 1; end
        16'b0101100011110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000010000000000000000000; ec = 1; end
        16'b1000011000100111:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000000100000000000000000000; ec = 1; end
        16'b1011011001101010:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000001000000000000000000000; ec = 1; end
        16'b1101011011110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000010000000000000000000000; ec = 1; end
        16'b0001011111000100:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000000100000000000000000000000; ec = 1; end
        16'b0001100001000001:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000001000000000000000000000000; ec = 1; end
        16'b0000011101001011:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000010000000000000000000000000; ec = 1; end
        16'b0011100101011111:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000000100000000000000000000000000; ec = 1; end
        16'b0100010101110111:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000001000000000000000000000000000; ec = 1; end
        16'b1011110100100111:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000010000000000000000000000000000; ec = 1; end
        16'b1100000001101010:begin data = code ^ 80'b00000000000000000000000000000000000000000000010000100000000000000000000000000000; ec = 1; end
        16'b0011101011110000:begin data = code ^ 80'b00000000000000000000000000000000000000000000010001000000000000000000000000000000; ec = 1; end
        16'b0100001000101001:begin data = code ^ 80'b00000000000000000000000000000000000000000000010010000000000000000000000000000000; ec = 1; end
        16'b1011001110011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000010100000000000000000000000000000000; ec = 1; end
        16'b1101110100010010:begin data = code ^ 80'b00000000000000000000000000000000000000000000011000000000000000000000000000000000; ec = 1; end
        16'b1010000111010100:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000000001; ec = 1; end
        16'b1010000111010111:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000000010; ec = 1; end
        16'b1010000111010001:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000000100; ec = 1; end
        16'b1010000111011101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000001000; ec = 1; end
        16'b1010000111000101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000010000; ec = 1; end
        16'b1010000111110101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000000100000; ec = 1; end
        16'b1010000110010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000001000000; ec = 1; end
        16'b1010000101010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000010000000; ec = 1; end
        16'b1010000011010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000000100000000; ec = 1; end
        16'b1010001111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000001000000000; ec = 1; end
        16'b1010010111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000010000000000; ec = 1; end
        16'b1010100111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000000100000000000; ec = 1; end
        16'b1011000111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000001000000000000; ec = 1; end
        16'b1000000111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000010000000000000; ec = 1; end
        16'b1110000111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000000100000000000000; ec = 1; end
        16'b0010000111010101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000001000000000000000; ec = 1; end
        16'b0010110000111000:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000010000000000000000; ec = 1; end
        16'b0011011111100010:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000000100000000000000000; ec = 1; end
        16'b0000000001010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000001000000000000000000; ec = 1; end
        16'b0110111100111110:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000010000000000000000000; ec = 1; end
        16'b1011000111101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000000100000000000000000000; ec = 1; end
        16'b1000000110100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000001000000000000000000000; ec = 1; end
        16'b1110000100111001:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000010000000000000000000000; ec = 1; end
        16'b0010000000001101:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000000100000000000000000000000; ec = 1; end
        16'b0010111110001000:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000001000000000000000000000000; ec = 1; end
        16'b0011000010000010:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000010000000000000000000000000; ec = 1; end
        16'b0000111010010110:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000000100000000000000000000000000; ec = 1; end
        16'b0111001010111110:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000001000000000000000000000000000; ec = 1; end
        16'b1000101011101110:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000010000000000000000000000000000; ec = 1; end
        16'b1111011110100011:begin data = code ^ 80'b00000000000000000000000000000000000000000000100000100000000000000000000000000000; ec = 1; end
        16'b0000110100111001:begin data = code ^ 80'b00000000000000000000000000000000000000000000100001000000000000000000000000000000; ec = 1; end
        16'b0111010111100000:begin data = code ^ 80'b00000000000000000000000000000000000000000000100010000000000000000000000000000000; ec = 1; end
        16'b1000010001010010:begin data = code ^ 80'b00000000000000000000000000000000000000000000100100000000000000000000000000000000; ec = 1; end
        16'b1110101011011011:begin data = code ^ 80'b00000000000000000000000000000000000000000000101000000000000000000000000000000000; ec = 1; end
        16'b0011011111001001:begin data = code ^ 80'b00000000000000000000000000000000000000000000110000000000000000000000000000000000; ec = 1; end
        16'b1100111001000110:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000000001; ec = 1; end
        16'b1100111001000101:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000000010; ec = 1; end
        16'b1100111001000011:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000000100; ec = 1; end
        16'b1100111001001111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000001000; ec = 1; end
        16'b1100111001010111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000010000; ec = 1; end
        16'b1100111001100111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000000100000; ec = 1; end
        16'b1100111000000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000001000000; ec = 1; end
        16'b1100111011000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000010000000; ec = 1; end
        16'b1100111101000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000000100000000; ec = 1; end
        16'b1100110001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000001000000000; ec = 1; end
        16'b1100101001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000010000000000; ec = 1; end
        16'b1100011001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000000100000000000; ec = 1; end
        16'b1101111001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000001000000000000; ec = 1; end
        16'b1110111001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000010000000000000; ec = 1; end
        16'b1000111001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000000100000000000000; ec = 1; end
        16'b0100111001000111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000001000000000000000; ec = 1; end
        16'b0100001110101010:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000010000000000000000; ec = 1; end
        16'b0101100001110000:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000000100000000000000000; ec = 1; end
        16'b0110111111000100:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000001000000000000000000; ec = 1; end
        16'b0000000010101100:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000010000000000000000000; ec = 1; end
        16'b1101111001111100:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000000100000000000000000000; ec = 1; end
        16'b1110111000110001:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000001000000000000000000000; ec = 1; end
        16'b1000111010101011:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000010000000000000000000000; ec = 1; end
        16'b0100111110011111:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000000100000000000000000000000; ec = 1; end
        16'b0100000000011010:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000001000000000000000000000000; ec = 1; end
        16'b0101111100010000:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000010000000000000000000000000; ec = 1; end
        16'b0110000100000100:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000000100000000000000000000000000; ec = 1; end
        16'b0001110100101100:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000001000000000000000000000000000; ec = 1; end
        16'b1110010101111100:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000010000000000000000000000000000; ec = 1; end
        16'b1001100000110001:begin data = code ^ 80'b00000000000000000000000000000000000000000001000000100000000000000000000000000000; ec = 1; end
        16'b0110001010101011:begin data = code ^ 80'b00000000000000000000000000000000000000000001000001000000000000000000000000000000; ec = 1; end
        16'b0001101001110010:begin data = code ^ 80'b00000000000000000000000000000000000000000001000010000000000000000000000000000000; ec = 1; end
        16'b1110101111000000:begin data = code ^ 80'b00000000000000000000000000000000000000000001000100000000000000000000000000000000; ec = 1; end
        16'b1000010101001001:begin data = code ^ 80'b00000000000000000000000000000000000000000001001000000000000000000000000000000000; ec = 1; end
        16'b0101100001011011:begin data = code ^ 80'b00000000000000000000000000000000000000000001010000000000000000000000000000000000; ec = 1; end
        16'b0110111110010010:begin data = code ^ 80'b00000000000000000000000000000000000000000001100000000000000000000000000000000000; ec = 1; end
        16'b0001000101100010:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000000001; ec = 1; end
        16'b0001000101100001:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000000010; ec = 1; end
        16'b0001000101100111:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000000100; ec = 1; end
        16'b0001000101101011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000001000; ec = 1; end
        16'b0001000101110011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000010000; ec = 1; end
        16'b0001000101000011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000000100000; ec = 1; end
        16'b0001000100100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000001000000; ec = 1; end
        16'b0001000111100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000010000000; ec = 1; end
        16'b0001000001100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000000100000000; ec = 1; end
        16'b0001001101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000001000000000; ec = 1; end
        16'b0001010101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000010000000000; ec = 1; end
        16'b0001100101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000000100000000000; ec = 1; end
        16'b0000000101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000001000000000000; ec = 1; end
        16'b0011000101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000010000000000000; ec = 1; end
        16'b0101000101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000000100000000000000; ec = 1; end
        16'b1001000101100011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000001000000000000000; ec = 1; end
        16'b1001110010001110:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000010000000000000000; ec = 1; end
        16'b1000011101010100:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000000100000000000000000; ec = 1; end
        16'b1011000011100000:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000001000000000000000000; ec = 1; end
        16'b1101111110001000:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000010000000000000000000; ec = 1; end
        16'b0000000101011000:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000000100000000000000000000; ec = 1; end
        16'b0011000100010101:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000001000000000000000000000; ec = 1; end
        16'b0101000110001111:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000010000000000000000000000; ec = 1; end
        16'b1001000010111011:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000000100000000000000000000000; ec = 1; end
        16'b1001111100111110:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000001000000000000000000000000; ec = 1; end
        16'b1000000000110100:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000010000000000000000000000000; ec = 1; end
        16'b1011111000100000:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000000100000000000000000000000000; ec = 1; end
        16'b1100001000001000:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000001000000000000000000000000000; ec = 1; end
        16'b0011101001011000:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000010000000000000000000000000000; ec = 1; end
        16'b0100011100010101:begin data = code ^ 80'b00000000000000000000000000000000000000000010000000100000000000000000000000000000; ec = 1; end
        16'b1011110110001111:begin data = code ^ 80'b00000000000000000000000000000000000000000010000001000000000000000000000000000000; ec = 1; end
        16'b1100010101010110:begin data = code ^ 80'b00000000000000000000000000000000000000000010000010000000000000000000000000000000; ec = 1; end
        16'b0011010011100100:begin data = code ^ 80'b00000000000000000000000000000000000000000010000100000000000000000000000000000000; ec = 1; end
        16'b0101101001101101:begin data = code ^ 80'b00000000000000000000000000000000000000000010001000000000000000000000000000000000; ec = 1; end
        16'b1000011101111111:begin data = code ^ 80'b00000000000000000000000000000000000000000010010000000000000000000000000000000000; ec = 1; end
        16'b1011000010110110:begin data = code ^ 80'b00000000000000000000000000000000000000000010100000000000000000000000000000000000; ec = 1; end
        16'b1101111100100100:begin data = code ^ 80'b00000000000000000000000000000000000000000011000000000000000000000000000000000000; ec = 1; end
        16'b0010001011000111:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000000001; ec = 1; end
        16'b0010001011000100:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000000010; ec = 1; end
        16'b0010001011000010:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000000100; ec = 1; end
        16'b0010001011001110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000001000; ec = 1; end
        16'b0010001011010110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000010000; ec = 1; end
        16'b0010001011100110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000000100000; ec = 1; end
        16'b0010001010000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000001000000; ec = 1; end
        16'b0010001001000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000010000000; ec = 1; end
        16'b0010001111000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000000100000000; ec = 1; end
        16'b0010000011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000001000000000; ec = 1; end
        16'b0010011011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000010000000000; ec = 1; end
        16'b0010101011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000000100000000000; ec = 1; end
        16'b0011001011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000001000000000000; ec = 1; end
        16'b0000001011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000010000000000000; ec = 1; end
        16'b0110001011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000000100000000000000; ec = 1; end
        16'b1010001011000110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000001000000000000000; ec = 1; end
        16'b1010111100101011:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000010000000000000000; ec = 1; end
        16'b1011010011110001:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000000100000000000000000; ec = 1; end
        16'b1000001101000101:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000001000000000000000000; ec = 1; end
        16'b1110110000101101:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000010000000000000000000; ec = 1; end
        16'b0011001011111101:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000000100000000000000000000; ec = 1; end
        16'b0000001010110000:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000001000000000000000000000; ec = 1; end
        16'b0110001000101010:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000010000000000000000000000; ec = 1; end
        16'b1010001100011110:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000000100000000000000000000000; ec = 1; end
        16'b1010110010011011:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000001000000000000000000000000; ec = 1; end
        16'b1011001110010001:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000010000000000000000000000000; ec = 1; end
        16'b1000110110000101:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000000100000000000000000000000000; ec = 1; end
        16'b1111000110101101:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000001000000000000000000000000000; ec = 1; end
        16'b0000100111111101:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000010000000000000000000000000000; ec = 1; end
        16'b0111010010110000:begin data = code ^ 80'b00000000000000000000000000000000000000000100000000100000000000000000000000000000; ec = 1; end
        16'b1000111000101010:begin data = code ^ 80'b00000000000000000000000000000000000000000100000001000000000000000000000000000000; ec = 1; end
        16'b1111011011110011:begin data = code ^ 80'b00000000000000000000000000000000000000000100000010000000000000000000000000000000; ec = 1; end
        16'b0000011101000001:begin data = code ^ 80'b00000000000000000000000000000000000000000100000100000000000000000000000000000000; ec = 1; end
        16'b0110100111001000:begin data = code ^ 80'b00000000000000000000000000000000000000000100001000000000000000000000000000000000; ec = 1; end
        16'b1011010011011010:begin data = code ^ 80'b00000000000000000000000000000000000000000100010000000000000000000000000000000000; ec = 1; end
        16'b1000001100010011:begin data = code ^ 80'b00000000000000000000000000000000000000000100100000000000000000000000000000000000; ec = 1; end
        16'b1110110010000001:begin data = code ^ 80'b00000000000000000000000000000000000000000101000000000000000000000000000000000000; ec = 1; end
        16'b0011001110100101:begin data = code ^ 80'b00000000000000000000000000000000000000000110000000000000000000000000000000000000; ec = 1; end
        16'b0100010110001101:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000000001; ec = 1; end
        16'b0100010110001110:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000000010; ec = 1; end
        16'b0100010110001000:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000000100; ec = 1; end
        16'b0100010110000100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000001000; ec = 1; end
        16'b0100010110011100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000010000; ec = 1; end
        16'b0100010110101100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000000100000; ec = 1; end
        16'b0100010111001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000001000000; ec = 1; end
        16'b0100010100001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000010000000; ec = 1; end
        16'b0100010010001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000000100000000; ec = 1; end
        16'b0100011110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000001000000000; ec = 1; end
        16'b0100000110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000010000000000; ec = 1; end
        16'b0100110110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000000100000000000; ec = 1; end
        16'b0101010110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000001000000000000; ec = 1; end
        16'b0110010110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000010000000000000; ec = 1; end
        16'b0000010110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000000100000000000000; ec = 1; end
        16'b1100010110001100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000001000000000000000; ec = 1; end
        16'b1100100001100001:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000010000000000000000; ec = 1; end
        16'b1101001110111011:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000000100000000000000000; ec = 1; end
        16'b1110010000001111:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000001000000000000000000; ec = 1; end
        16'b1000101101100111:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000010000000000000000000; ec = 1; end
        16'b0101010110110111:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000000100000000000000000000; ec = 1; end
        16'b0110010111111010:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000001000000000000000000000; ec = 1; end
        16'b0000010101100000:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000010000000000000000000000; ec = 1; end
        16'b1100010001010100:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000000100000000000000000000000; ec = 1; end
        16'b1100101111010001:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000001000000000000000000000000; ec = 1; end
        16'b1101010011011011:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000010000000000000000000000000; ec = 1; end
        16'b1110101011001111:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000000100000000000000000000000000; ec = 1; end
        16'b1001011011100111:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000001000000000000000000000000000; ec = 1; end
        16'b0110111010110111:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000010000000000000000000000000000; ec = 1; end
        16'b0001001111111010:begin data = code ^ 80'b00000000000000000000000000000000000000001000000000100000000000000000000000000000; ec = 1; end
        16'b1110100101100000:begin data = code ^ 80'b00000000000000000000000000000000000000001000000001000000000000000000000000000000; ec = 1; end
        16'b1001000110111001:begin data = code ^ 80'b00000000000000000000000000000000000000001000000010000000000000000000000000000000; ec = 1; end
        16'b0110000000001011:begin data = code ^ 80'b00000000000000000000000000000000000000001000000100000000000000000000000000000000; ec = 1; end
        16'b0000111010000010:begin data = code ^ 80'b00000000000000000000000000000000000000001000001000000000000000000000000000000000; ec = 1; end
        16'b1101001110010000:begin data = code ^ 80'b00000000000000000000000000000000000000001000010000000000000000000000000000000000; ec = 1; end
        16'b1110010001011001:begin data = code ^ 80'b00000000000000000000000000000000000000001000100000000000000000000000000000000000; ec = 1; end
        16'b1000101111001011:begin data = code ^ 80'b00000000000000000000000000000000000000001001000000000000000000000000000000000000; ec = 1; end
        16'b0101010011101111:begin data = code ^ 80'b00000000000000000000000000000000000000001010000000000000000000000000000000000000; ec = 1; end
        16'b0110011101001010:begin data = code ^ 80'b00000000000000000000000000000000000000001100000000000000000000000000000000000000; ec = 1; end
        16'b1000101100011001:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000000001; ec = 1; end
        16'b1000101100011010:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000000010; ec = 1; end
        16'b1000101100011100:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000000100; ec = 1; end
        16'b1000101100010000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000001000; ec = 1; end
        16'b1000101100001000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000010000; ec = 1; end
        16'b1000101100111000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000000100000; ec = 1; end
        16'b1000101101011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000001000000; ec = 1; end
        16'b1000101110011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000010000000; ec = 1; end
        16'b1000101000011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000000100000000; ec = 1; end
        16'b1000100100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000001000000000; ec = 1; end
        16'b1000111100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000010000000000; ec = 1; end
        16'b1000001100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000000100000000000; ec = 1; end
        16'b1001101100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000001000000000000; ec = 1; end
        16'b1010101100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000010000000000000; ec = 1; end
        16'b1100101100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000000100000000000000; ec = 1; end
        16'b0000101100011000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000001000000000000000; ec = 1; end
        16'b0000011011110101:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000010000000000000000; ec = 1; end
        16'b0001110100101111:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000000100000000000000000; ec = 1; end
        16'b0010101010011011:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000001000000000000000000; ec = 1; end
        16'b0100010111110011:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000010000000000000000000; ec = 1; end
        16'b1001101100100011:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000000100000000000000000000; ec = 1; end
        16'b1010101101101110:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000001000000000000000000000; ec = 1; end
        16'b1100101111110100:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000010000000000000000000000; ec = 1; end
        16'b0000101011000000:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000000100000000000000000000000; ec = 1; end
        16'b0000010101000101:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000001000000000000000000000000; ec = 1; end
        16'b0001101001001111:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000010000000000000000000000000; ec = 1; end
        16'b0010010001011011:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000000100000000000000000000000000; ec = 1; end
        16'b0101100001110011:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000001000000000000000000000000000; ec = 1; end
        16'b1010000000100011:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000010000000000000000000000000000; ec = 1; end
        16'b1101110101101110:begin data = code ^ 80'b00000000000000000000000000000000000000010000000000100000000000000000000000000000; ec = 1; end
        16'b0010011111110100:begin data = code ^ 80'b00000000000000000000000000000000000000010000000001000000000000000000000000000000; ec = 1; end
        16'b0101111100101101:begin data = code ^ 80'b00000000000000000000000000000000000000010000000010000000000000000000000000000000; ec = 1; end
        16'b1010111010011111:begin data = code ^ 80'b00000000000000000000000000000000000000010000000100000000000000000000000000000000; ec = 1; end
        16'b1100000000010110:begin data = code ^ 80'b00000000000000000000000000000000000000010000001000000000000000000000000000000000; ec = 1; end
        16'b0001110100000100:begin data = code ^ 80'b00000000000000000000000000000000000000010000010000000000000000000000000000000000; ec = 1; end
        16'b0010101011001101:begin data = code ^ 80'b00000000000000000000000000000000000000010000100000000000000000000000000000000000; ec = 1; end
        16'b0100010101011111:begin data = code ^ 80'b00000000000000000000000000000000000000010001000000000000000000000000000000000000; ec = 1; end
        16'b1001101001111011:begin data = code ^ 80'b00000000000000000000000000000000000000010010000000000000000000000000000000000000; ec = 1; end
        16'b1010100111011110:begin data = code ^ 80'b00000000000000000000000000000000000000010100000000000000000000000000000000000000; ec = 1; end
        16'b1100111010010100:begin data = code ^ 80'b00000000000000000000000000000000000000011000000000000000000000000000000000000000; ec = 1; end
        16'b1001101111011100:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000000001; ec = 1; end
        16'b1001101111011111:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000000010; ec = 1; end
        16'b1001101111011001:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000000100; ec = 1; end
        16'b1001101111010101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000001000; ec = 1; end
        16'b1001101111001101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000010000; ec = 1; end
        16'b1001101111111101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000000100000; ec = 1; end
        16'b1001101110011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000001000000; ec = 1; end
        16'b1001101101011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000010000000; ec = 1; end
        16'b1001101011011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000000100000000; ec = 1; end
        16'b1001100111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000001000000000; ec = 1; end
        16'b1001111111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000010000000000; ec = 1; end
        16'b1001001111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000000100000000000; ec = 1; end
        16'b1000101111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000001000000000000; ec = 1; end
        16'b1011101111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000010000000000000; ec = 1; end
        16'b1101101111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000000100000000000000; ec = 1; end
        16'b0001101111011101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000001000000000000000; ec = 1; end
        16'b0001011000110000:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000010000000000000000; ec = 1; end
        16'b0000110111101010:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000000100000000000000000; ec = 1; end
        16'b0011101001011110:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000001000000000000000000; ec = 1; end
        16'b0101010100110110:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000010000000000000000000; ec = 1; end
        16'b1000101111100110:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000000100000000000000000000; ec = 1; end
        16'b1011101110101011:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000001000000000000000000000; ec = 1; end
        16'b1101101100110001:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000010000000000000000000000; ec = 1; end
        16'b0001101000000101:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000000100000000000000000000000; ec = 1; end
        16'b0001010110000000:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000001000000000000000000000000; ec = 1; end
        16'b0000101010001010:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000010000000000000000000000000; ec = 1; end
        16'b0011010010011110:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000000100000000000000000000000000; ec = 1; end
        16'b0100100010110110:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000001000000000000000000000000000; ec = 1; end
        16'b1011000011100110:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000010000000000000000000000000000; ec = 1; end
        16'b1100110110101011:begin data = code ^ 80'b00000000000000000000000000000000000000100000000000100000000000000000000000000000; ec = 1; end
        16'b0011011100110001:begin data = code ^ 80'b00000000000000000000000000000000000000100000000001000000000000000000000000000000; ec = 1; end
        16'b0100111111101000:begin data = code ^ 80'b00000000000000000000000000000000000000100000000010000000000000000000000000000000; ec = 1; end
        16'b1011111001011010:begin data = code ^ 80'b00000000000000000000000000000000000000100000000100000000000000000000000000000000; ec = 1; end
        16'b1101000011010011:begin data = code ^ 80'b00000000000000000000000000000000000000100000001000000000000000000000000000000000; ec = 1; end
        16'b0000110111000001:begin data = code ^ 80'b00000000000000000000000000000000000000100000010000000000000000000000000000000000; ec = 1; end
        16'b0011101000001000:begin data = code ^ 80'b00000000000000000000000000000000000000100000100000000000000000000000000000000000; ec = 1; end
        16'b0101010110011010:begin data = code ^ 80'b00000000000000000000000000000000000000100001000000000000000000000000000000000000; ec = 1; end
        16'b1000101010111110:begin data = code ^ 80'b00000000000000000000000000000000000000100010000000000000000000000000000000000000; ec = 1; end
        16'b1011100100011011:begin data = code ^ 80'b00000000000000000000000000000000000000100100000000000000000000000000000000000000; ec = 1; end
        16'b1101111001010001:begin data = code ^ 80'b00000000000000000000000000000000000000101000000000000000000000000000000000000000; ec = 1; end
        16'b0001000011000101:begin data = code ^ 80'b00000000000000000000000000000000000000110000000000000000000000000000000000000000; ec = 1; end
        16'b1011101001010110:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000000001; ec = 1; end
        16'b1011101001010101:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000000010; ec = 1; end
        16'b1011101001010011:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000000100; ec = 1; end
        16'b1011101001011111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000001000; ec = 1; end
        16'b1011101001000111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000010000; ec = 1; end
        16'b1011101001110111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000000100000; ec = 1; end
        16'b1011101000010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000001000000; ec = 1; end
        16'b1011101011010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000010000000; ec = 1; end
        16'b1011101101010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000000100000000; ec = 1; end
        16'b1011100001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000001000000000; ec = 1; end
        16'b1011111001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000010000000000; ec = 1; end
        16'b1011001001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000000100000000000; ec = 1; end
        16'b1010101001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000001000000000000; ec = 1; end
        16'b1001101001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000010000000000000; ec = 1; end
        16'b1111101001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000000100000000000000; ec = 1; end
        16'b0011101001010111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000001000000000000000; ec = 1; end
        16'b0011011110111010:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000010000000000000000; ec = 1; end
        16'b0010110001100000:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000000100000000000000000; ec = 1; end
        16'b0001101111010100:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000001000000000000000000; ec = 1; end
        16'b0111010010111100:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000010000000000000000000; ec = 1; end
        16'b1010101001101100:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000000100000000000000000000; ec = 1; end
        16'b1001101000100001:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000001000000000000000000000; ec = 1; end
        16'b1111101010111011:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000010000000000000000000000; ec = 1; end
        16'b0011101110001111:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000000100000000000000000000000; ec = 1; end
        16'b0011010000001010:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000001000000000000000000000000; ec = 1; end
        16'b0010101100000000:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000010000000000000000000000000; ec = 1; end
        16'b0001010100010100:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000000100000000000000000000000000; ec = 1; end
        16'b0110100100111100:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000001000000000000000000000000000; ec = 1; end
        16'b1001000101101100:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000010000000000000000000000000000; ec = 1; end
        16'b1110110000100001:begin data = code ^ 80'b00000000000000000000000000000000000001000000000000100000000000000000000000000000; ec = 1; end
        16'b0001011010111011:begin data = code ^ 80'b00000000000000000000000000000000000001000000000001000000000000000000000000000000; ec = 1; end
        16'b0110111001100010:begin data = code ^ 80'b00000000000000000000000000000000000001000000000010000000000000000000000000000000; ec = 1; end
        16'b1001111111010000:begin data = code ^ 80'b00000000000000000000000000000000000001000000000100000000000000000000000000000000; ec = 1; end
        16'b1111000101011001:begin data = code ^ 80'b00000000000000000000000000000000000001000000001000000000000000000000000000000000; ec = 1; end
        16'b0010110001001011:begin data = code ^ 80'b00000000000000000000000000000000000001000000010000000000000000000000000000000000; ec = 1; end
        16'b0001101110000010:begin data = code ^ 80'b00000000000000000000000000000000000001000000100000000000000000000000000000000000; ec = 1; end
        16'b0111010000010000:begin data = code ^ 80'b00000000000000000000000000000000000001000001000000000000000000000000000000000000; ec = 1; end
        16'b1010101100110100:begin data = code ^ 80'b00000000000000000000000000000000000001000010000000000000000000000000000000000000; ec = 1; end
        16'b1001100010010001:begin data = code ^ 80'b00000000000000000000000000000000000001000100000000000000000000000000000000000000; ec = 1; end
        16'b1111111111011011:begin data = code ^ 80'b00000000000000000000000000000000000001001000000000000000000000000000000000000000; ec = 1; end
        16'b0011000101001111:begin data = code ^ 80'b00000000000000000000000000000000000001010000000000000000000000000000000000000000; ec = 1; end
        16'b0010000110001010:begin data = code ^ 80'b00000000000000000000000000000000000001100000000000000000000000000000000000000000; ec = 1; end
        16'b1111100101000010:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000000001; ec = 1; end
        16'b1111100101000001:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000000010; ec = 1; end
        16'b1111100101000111:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000000100; ec = 1; end
        16'b1111100101001011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000001000; ec = 1; end
        16'b1111100101010011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000010000; ec = 1; end
        16'b1111100101100011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000000100000; ec = 1; end
        16'b1111100100000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000001000000; ec = 1; end
        16'b1111100111000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000010000000; ec = 1; end
        16'b1111100001000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000000100000000; ec = 1; end
        16'b1111101101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000001000000000; ec = 1; end
        16'b1111110101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000010000000000; ec = 1; end
        16'b1111000101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000000100000000000; ec = 1; end
        16'b1110100101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000001000000000000; ec = 1; end
        16'b1101100101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000010000000000000; ec = 1; end
        16'b1011100101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000000100000000000000; ec = 1; end
        16'b0111100101000011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000001000000000000000; ec = 1; end
        16'b0111010010101110:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000010000000000000000; ec = 1; end
        16'b0110111101110100:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000000100000000000000000; ec = 1; end
        16'b0101100011000000:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000001000000000000000000; ec = 1; end
        16'b0011011110101000:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000010000000000000000000; ec = 1; end
        16'b1110100101111000:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000000100000000000000000000; ec = 1; end
        16'b1101100100110101:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000001000000000000000000000; ec = 1; end
        16'b1011100110101111:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000010000000000000000000000; ec = 1; end
        16'b0111100010011011:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000000100000000000000000000000; ec = 1; end
        16'b0111011100011110:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000001000000000000000000000000; ec = 1; end
        16'b0110100000010100:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000010000000000000000000000000; ec = 1; end
        16'b0101011000000000:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000000100000000000000000000000000; ec = 1; end
        16'b0010101000101000:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000001000000000000000000000000000; ec = 1; end
        16'b1101001001111000:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000010000000000000000000000000000; ec = 1; end
        16'b1010111100110101:begin data = code ^ 80'b00000000000000000000000000000000000010000000000000100000000000000000000000000000; ec = 1; end
        16'b0101010110101111:begin data = code ^ 80'b00000000000000000000000000000000000010000000000001000000000000000000000000000000; ec = 1; end
        16'b0010110101110110:begin data = code ^ 80'b00000000000000000000000000000000000010000000000010000000000000000000000000000000; ec = 1; end
        16'b1101110011000100:begin data = code ^ 80'b00000000000000000000000000000000000010000000000100000000000000000000000000000000; ec = 1; end
        16'b1011001001001101:begin data = code ^ 80'b00000000000000000000000000000000000010000000001000000000000000000000000000000000; ec = 1; end
        16'b0110111101011111:begin data = code ^ 80'b00000000000000000000000000000000000010000000010000000000000000000000000000000000; ec = 1; end
        16'b0101100010010110:begin data = code ^ 80'b00000000000000000000000000000000000010000000100000000000000000000000000000000000; ec = 1; end
        16'b0011011100000100:begin data = code ^ 80'b00000000000000000000000000000000000010000001000000000000000000000000000000000000; ec = 1; end
        16'b1110100000100000:begin data = code ^ 80'b00000000000000000000000000000000000010000010000000000000000000000000000000000000; ec = 1; end
        16'b1101101110000101:begin data = code ^ 80'b00000000000000000000000000000000000010000100000000000000000000000000000000000000; ec = 1; end
        16'b1011110011001111:begin data = code ^ 80'b00000000000000000000000000000000000010001000000000000000000000000000000000000000; ec = 1; end
        16'b0111001001011011:begin data = code ^ 80'b00000000000000000000000000000000000010010000000000000000000000000000000000000000; ec = 1; end
        16'b0110001010011110:begin data = code ^ 80'b00000000000000000000000000000000000010100000000000000000000000000000000000000000; ec = 1; end
        16'b0100001100010100:begin data = code ^ 80'b00000000000000000000000000000000000011000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111101101010:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000000001; ec = 1; end
        16'b0111111101101001:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000000010; ec = 1; end
        16'b0111111101101111:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000000100; ec = 1; end
        16'b0111111101100011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000001000; ec = 1; end
        16'b0111111101111011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000010000; ec = 1; end
        16'b0111111101001011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000000100000; ec = 1; end
        16'b0111111100101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000001000000; ec = 1; end
        16'b0111111111101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000010000000; ec = 1; end
        16'b0111111001101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000000100000000; ec = 1; end
        16'b0111110101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000001000000000; ec = 1; end
        16'b0111101101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000010000000000; ec = 1; end
        16'b0111011101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000000100000000000; ec = 1; end
        16'b0110111101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000001000000000000; ec = 1; end
        16'b0101111101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000010000000000000; ec = 1; end
        16'b0011111101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000000100000000000000; ec = 1; end
        16'b1111111101101011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000001000000000000000; ec = 1; end
        16'b1111001010000110:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000010000000000000000; ec = 1; end
        16'b1110100101011100:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000000100000000000000000; ec = 1; end
        16'b1101111011101000:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000001000000000000000000; ec = 1; end
        16'b1011000110000000:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000010000000000000000000; ec = 1; end
        16'b0110111101010000:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000000100000000000000000000; ec = 1; end
        16'b0101111100011101:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000001000000000000000000000; ec = 1; end
        16'b0011111110000111:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000010000000000000000000000; ec = 1; end
        16'b1111111010110011:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000000100000000000000000000000; ec = 1; end
        16'b1111000100110110:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000001000000000000000000000000; ec = 1; end
        16'b1110111000111100:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000010000000000000000000000000; ec = 1; end
        16'b1101000000101000:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000000100000000000000000000000000; ec = 1; end
        16'b1010110000000000:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000001000000000000000000000000000; ec = 1; end
        16'b0101010001010000:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000010000000000000000000000000000; ec = 1; end
        16'b0010100100011101:begin data = code ^ 80'b00000000000000000000000000000000000100000000000000100000000000000000000000000000; ec = 1; end
        16'b1101001110000111:begin data = code ^ 80'b00000000000000000000000000000000000100000000000001000000000000000000000000000000; ec = 1; end
        16'b1010101101011110:begin data = code ^ 80'b00000000000000000000000000000000000100000000000010000000000000000000000000000000; ec = 1; end
        16'b0101101011101100:begin data = code ^ 80'b00000000000000000000000000000000000100000000000100000000000000000000000000000000; ec = 1; end
        16'b0011010001100101:begin data = code ^ 80'b00000000000000000000000000000000000100000000001000000000000000000000000000000000; ec = 1; end
        16'b1110100101110111:begin data = code ^ 80'b00000000000000000000000000000000000100000000010000000000000000000000000000000000; ec = 1; end
        16'b1101111010111110:begin data = code ^ 80'b00000000000000000000000000000000000100000000100000000000000000000000000000000000; ec = 1; end
        16'b1011000100101100:begin data = code ^ 80'b00000000000000000000000000000000000100000001000000000000000000000000000000000000; ec = 1; end
        16'b0110111000001000:begin data = code ^ 80'b00000000000000000000000000000000000100000010000000000000000000000000000000000000; ec = 1; end
        16'b0101110110101101:begin data = code ^ 80'b00000000000000000000000000000000000100000100000000000000000000000000000000000000; ec = 1; end
        16'b0011101011100111:begin data = code ^ 80'b00000000000000000000000000000000000100001000000000000000000000000000000000000000; ec = 1; end
        16'b1111010001110011:begin data = code ^ 80'b00000000000000000000000000000000000100010000000000000000000000000000000000000000; ec = 1; end
        16'b1110010010110110:begin data = code ^ 80'b00000000000000000000000000000000000100100000000000000000000000000000000000000000; ec = 1; end
        16'b1100010100111100:begin data = code ^ 80'b00000000000000000000000000000000000101000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011000101000:begin data = code ^ 80'b00000000000000000000000000000000000110000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111011010111:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000000001; ec = 1; end
        16'b1111111011010100:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000000010; ec = 1; end
        16'b1111111011010010:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000000100; ec = 1; end
        16'b1111111011011110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000001000; ec = 1; end
        16'b1111111011000110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000010000; ec = 1; end
        16'b1111111011110110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000000100000; ec = 1; end
        16'b1111111010010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000001000000; ec = 1; end
        16'b1111111001010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000010000000; ec = 1; end
        16'b1111111111010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000000100000000; ec = 1; end
        16'b1111110011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000001000000000; ec = 1; end
        16'b1111101011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000010000000000; ec = 1; end
        16'b1111011011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000000100000000000; ec = 1; end
        16'b1110111011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000001000000000000; ec = 1; end
        16'b1101111011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000010000000000000; ec = 1; end
        16'b1011111011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000000100000000000000; ec = 1; end
        16'b0111111011010110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000001000000000000000; ec = 1; end
        16'b0111001100111011:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000010000000000000000; ec = 1; end
        16'b0110100011100001:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000000100000000000000000; ec = 1; end
        16'b0101111101010101:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000001000000000000000000; ec = 1; end
        16'b0011000000111101:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000010000000000000000000; ec = 1; end
        16'b1110111011101101:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000000100000000000000000000; ec = 1; end
        16'b1101111010100000:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000001000000000000000000000; ec = 1; end
        16'b1011111000111010:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000010000000000000000000000; ec = 1; end
        16'b0111111100001110:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000000100000000000000000000000; ec = 1; end
        16'b0111000010001011:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000001000000000000000000000000; ec = 1; end
        16'b0110111110000001:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000010000000000000000000000000; ec = 1; end
        16'b0101000110010101:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000000100000000000000000000000000; ec = 1; end
        16'b0010110110111101:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000001000000000000000000000000000; ec = 1; end
        16'b1101010111101101:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000010000000000000000000000000000; ec = 1; end
        16'b1010100010100000:begin data = code ^ 80'b00000000000000000000000000000000001000000000000000100000000000000000000000000000; ec = 1; end
        16'b0101001000111010:begin data = code ^ 80'b00000000000000000000000000000000001000000000000001000000000000000000000000000000; ec = 1; end
        16'b0010101011100011:begin data = code ^ 80'b00000000000000000000000000000000001000000000000010000000000000000000000000000000; ec = 1; end
        16'b1101101101010001:begin data = code ^ 80'b00000000000000000000000000000000001000000000000100000000000000000000000000000000; ec = 1; end
        16'b1011010111011000:begin data = code ^ 80'b00000000000000000000000000000000001000000000001000000000000000000000000000000000; ec = 1; end
        16'b0110100011001010:begin data = code ^ 80'b00000000000000000000000000000000001000000000010000000000000000000000000000000000; ec = 1; end
        16'b0101111100000011:begin data = code ^ 80'b00000000000000000000000000000000001000000000100000000000000000000000000000000000; ec = 1; end
        16'b0011000010010001:begin data = code ^ 80'b00000000000000000000000000000000001000000001000000000000000000000000000000000000; ec = 1; end
        16'b1110111110110101:begin data = code ^ 80'b00000000000000000000000000000000001000000010000000000000000000000000000000000000; ec = 1; end
        16'b1101110000010000:begin data = code ^ 80'b00000000000000000000000000000000001000000100000000000000000000000000000000000000; ec = 1; end
        16'b1011101101011010:begin data = code ^ 80'b00000000000000000000000000000000001000001000000000000000000000000000000000000000; ec = 1; end
        16'b0111010111001110:begin data = code ^ 80'b00000000000000000000000000000000001000010000000000000000000000000000000000000000; ec = 1; end
        16'b0110010100001011:begin data = code ^ 80'b00000000000000000000000000000000001000100000000000000000000000000000000000000000; ec = 1; end
        16'b0100010010000001:begin data = code ^ 80'b00000000000000000000000000000000001001000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011110010101:begin data = code ^ 80'b00000000000000000000000000000000001010000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000110111101:begin data = code ^ 80'b00000000000000000000000000000000001100000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000001000000:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000000001; ec = 1; end
        16'b0111000001000011:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000000010; ec = 1; end
        16'b0111000001000101:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000000100; ec = 1; end
        16'b0111000001001001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000001000; ec = 1; end
        16'b0111000001010001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000010000; ec = 1; end
        16'b0111000001100001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000000100000; ec = 1; end
        16'b0111000000000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000001000000; ec = 1; end
        16'b0111000011000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000010000000; ec = 1; end
        16'b0111000101000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000000100000000; ec = 1; end
        16'b0111001001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000001000000000; ec = 1; end
        16'b0111010001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000010000000000; ec = 1; end
        16'b0111100001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000000100000000000; ec = 1; end
        16'b0110000001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000001000000000000; ec = 1; end
        16'b0101000001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000010000000000000; ec = 1; end
        16'b0011000001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000000100000000000000; ec = 1; end
        16'b1111000001000001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000001000000000000000; ec = 1; end
        16'b1111110110101100:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000010000000000000000; ec = 1; end
        16'b1110011001110110:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000000100000000000000000; ec = 1; end
        16'b1101000111000010:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000001000000000000000000; ec = 1; end
        16'b1011111010101010:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000010000000000000000000; ec = 1; end
        16'b0110000001111010:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000000100000000000000000000; ec = 1; end
        16'b0101000000110111:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000001000000000000000000000; ec = 1; end
        16'b0011000010101101:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000010000000000000000000000; ec = 1; end
        16'b1111000110011001:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000000100000000000000000000000; ec = 1; end
        16'b1111111000011100:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000001000000000000000000000000; ec = 1; end
        16'b1110000100010110:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000010000000000000000000000000; ec = 1; end
        16'b1101111100000010:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000000100000000000000000000000000; ec = 1; end
        16'b1010001100101010:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000001000000000000000000000000000; ec = 1; end
        16'b0101101101111010:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000010000000000000000000000000000; ec = 1; end
        16'b0010011000110111:begin data = code ^ 80'b00000000000000000000000000000000010000000000000000100000000000000000000000000000; ec = 1; end
        16'b1101110010101101:begin data = code ^ 80'b00000000000000000000000000000000010000000000000001000000000000000000000000000000; ec = 1; end
        16'b1010010001110100:begin data = code ^ 80'b00000000000000000000000000000000010000000000000010000000000000000000000000000000; ec = 1; end
        16'b0101010111000110:begin data = code ^ 80'b00000000000000000000000000000000010000000000000100000000000000000000000000000000; ec = 1; end
        16'b0011101101001111:begin data = code ^ 80'b00000000000000000000000000000000010000000000001000000000000000000000000000000000; ec = 1; end
        16'b1110011001011101:begin data = code ^ 80'b00000000000000000000000000000000010000000000010000000000000000000000000000000000; ec = 1; end
        16'b1101000110010100:begin data = code ^ 80'b00000000000000000000000000000000010000000000100000000000000000000000000000000000; ec = 1; end
        16'b1011111000000110:begin data = code ^ 80'b00000000000000000000000000000000010000000001000000000000000000000000000000000000; ec = 1; end
        16'b0110000100100010:begin data = code ^ 80'b00000000000000000000000000000000010000000010000000000000000000000000000000000000; ec = 1; end
        16'b0101001010000111:begin data = code ^ 80'b00000000000000000000000000000000010000000100000000000000000000000000000000000000; ec = 1; end
        16'b0011010111001101:begin data = code ^ 80'b00000000000000000000000000000000010000001000000000000000000000000000000000000000; ec = 1; end
        16'b1111101101011001:begin data = code ^ 80'b00000000000000000000000000000000010000010000000000000000000000000000000000000000; ec = 1; end
        16'b1110101110011100:begin data = code ^ 80'b00000000000000000000000000000000010000100000000000000000000000000000000000000000; ec = 1; end
        16'b1100101000010110:begin data = code ^ 80'b00000000000000000000000000000000010001000000000000000000000000000000000000000000; ec = 1; end
        16'b1000100100000010:begin data = code ^ 80'b00000000000000000000000000000000010010000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111100101010:begin data = code ^ 80'b00000000000000000000000000000000010100000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111010010111:begin data = code ^ 80'b00000000000000000000000000000000011000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000010000011:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000000001; ec = 1; end
        16'b1110000010000000:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000000010; ec = 1; end
        16'b1110000010000110:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000000100; ec = 1; end
        16'b1110000010001010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000001000; ec = 1; end
        16'b1110000010010010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000010000; ec = 1; end
        16'b1110000010100010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000000100000; ec = 1; end
        16'b1110000011000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000001000000; ec = 1; end
        16'b1110000000000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000010000000; ec = 1; end
        16'b1110000110000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000000100000000; ec = 1; end
        16'b1110001010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000001000000000; ec = 1; end
        16'b1110010010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000010000000000; ec = 1; end
        16'b1110100010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000000100000000000; ec = 1; end
        16'b1111000010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000001000000000000; ec = 1; end
        16'b1100000010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000010000000000000; ec = 1; end
        16'b1010000010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000000100000000000000; ec = 1; end
        16'b0110000010000010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000001000000000000000; ec = 1; end
        16'b0110110101101111:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000010000000000000000; ec = 1; end
        16'b0111011010110101:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000000100000000000000000; ec = 1; end
        16'b0100000100000001:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000001000000000000000000; ec = 1; end
        16'b0010111001101001:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000010000000000000000000; ec = 1; end
        16'b1111000010111001:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000000100000000000000000000; ec = 1; end
        16'b1100000011110100:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000001000000000000000000000; ec = 1; end
        16'b1010000001101110:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000010000000000000000000000; ec = 1; end
        16'b0110000101011010:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000000100000000000000000000000; ec = 1; end
        16'b0110111011011111:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000001000000000000000000000000; ec = 1; end
        16'b0111000111010101:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000010000000000000000000000000; ec = 1; end
        16'b0100111111000001:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000000100000000000000000000000000; ec = 1; end
        16'b0011001111101001:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000001000000000000000000000000000; ec = 1; end
        16'b1100101110111001:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000010000000000000000000000000000; ec = 1; end
        16'b1011011011110100:begin data = code ^ 80'b00000000000000000000000000000000100000000000000000100000000000000000000000000000; ec = 1; end
        16'b0100110001101110:begin data = code ^ 80'b00000000000000000000000000000000100000000000000001000000000000000000000000000000; ec = 1; end
        16'b0011010010110111:begin data = code ^ 80'b00000000000000000000000000000000100000000000000010000000000000000000000000000000; ec = 1; end
        16'b1100010100000101:begin data = code ^ 80'b00000000000000000000000000000000100000000000000100000000000000000000000000000000; ec = 1; end
        16'b1010101110001100:begin data = code ^ 80'b00000000000000000000000000000000100000000000001000000000000000000000000000000000; ec = 1; end
        16'b0111011010011110:begin data = code ^ 80'b00000000000000000000000000000000100000000000010000000000000000000000000000000000; ec = 1; end
        16'b0100000101010111:begin data = code ^ 80'b00000000000000000000000000000000100000000000100000000000000000000000000000000000; ec = 1; end
        16'b0010111011000101:begin data = code ^ 80'b00000000000000000000000000000000100000000001000000000000000000000000000000000000; ec = 1; end
        16'b1111000111100001:begin data = code ^ 80'b00000000000000000000000000000000100000000010000000000000000000000000000000000000; ec = 1; end
        16'b1100001001000100:begin data = code ^ 80'b00000000000000000000000000000000100000000100000000000000000000000000000000000000; ec = 1; end
        16'b1010010100001110:begin data = code ^ 80'b00000000000000000000000000000000100000001000000000000000000000000000000000000000; ec = 1; end
        16'b0110101110011010:begin data = code ^ 80'b00000000000000000000000000000000100000010000000000000000000000000000000000000000; ec = 1; end
        16'b0111101101011111:begin data = code ^ 80'b00000000000000000000000000000000100000100000000000000000000000000000000000000000; ec = 1; end
        16'b0101101011010101:begin data = code ^ 80'b00000000000000000000000000000000100001000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100111000001:begin data = code ^ 80'b00000000000000000000000000000000100010000000000000000000000000000000000000000000; ec = 1; end
        16'b1001111111101001:begin data = code ^ 80'b00000000000000000000000000000000100100000000000000000000000000000000000000000000; ec = 1; end
        16'b0001111001010100:begin data = code ^ 80'b00000000000000000000000000000000101000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000011000011:begin data = code ^ 80'b00000000000000000000000000000000110000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110011101000:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0100110011101011:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0100110011101101:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0100110011100001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0100110011111001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0100110011001001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0100110010101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0100110001101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0100110111101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0100111011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0100100011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0100010011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0101110011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0110110011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0000110011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1100110011101001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1100000100000100:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1101101011011110:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1110110101101010:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1000001000000010:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0101110011010010:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0110110010011111:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0000110000000101:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1100110100110001:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1100001010110100:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1101110110111110:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1110001110101010:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1001111110000010:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0110011111010010:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0001101010011111:begin data = code ^ 80'b00000000000000000000000000000001000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1110000000000101:begin data = code ^ 80'b00000000000000000000000000000001000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1001100011011100:begin data = code ^ 80'b00000000000000000000000000000001000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0110100101101110:begin data = code ^ 80'b00000000000000000000000000000001000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0000011111100111:begin data = code ^ 80'b00000000000000000000000000000001000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1101101011110101:begin data = code ^ 80'b00000000000000000000000000000001000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1110110100111100:begin data = code ^ 80'b00000000000000000000000000000001000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1000001010101110:begin data = code ^ 80'b00000000000000000000000000000001000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0101110110001010:begin data = code ^ 80'b00000000000000000000000000000001000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0110111000101111:begin data = code ^ 80'b00000000000000000000000000000001000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0000100101100101:begin data = code ^ 80'b00000000000000000000000000000001000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1100011111110001:begin data = code ^ 80'b00000000000000000000000000000001000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1101011100110100:begin data = code ^ 80'b00000000000000000000000000000001000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1111011010111110:begin data = code ^ 80'b00000000000000000000000000000001000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1011010110101010:begin data = code ^ 80'b00000000000000000000000000000001000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001110000010:begin data = code ^ 80'b00000000000000000000000000000001000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1011001000111111:begin data = code ^ 80'b00000000000000000000000000000001001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011110010101000:begin data = code ^ 80'b00000000000000000000000000000001010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010110001101011:begin data = code ^ 80'b00000000000000000000000000000001100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100111010011:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1001100111010000:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1001100111010110:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1001100111011010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1001100111000010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1001100111110010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1001100110010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1001100101010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1001100011010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1001101111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1001110111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1001000111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1000100111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1011100111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1101100111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0001100111010010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0001010000111111:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0000111111100101:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0011100001010001:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0101011100111001:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1000100111101001:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1011100110100100:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1101100100111110:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0001100000001010:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0001011110001111:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0000100010000101:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0011011010010001:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0100101010111001:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1011001011101001:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1100111110100100:begin data = code ^ 80'b00000000000000000000000000000010000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0011010100111110:begin data = code ^ 80'b00000000000000000000000000000010000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0100110111100111:begin data = code ^ 80'b00000000000000000000000000000010000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1011110001010101:begin data = code ^ 80'b00000000000000000000000000000010000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1101001011011100:begin data = code ^ 80'b00000000000000000000000000000010000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0000111111001110:begin data = code ^ 80'b00000000000000000000000000000010000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0011100000000111:begin data = code ^ 80'b00000000000000000000000000000010000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0101011110010101:begin data = code ^ 80'b00000000000000000000000000000010000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1000100010110001:begin data = code ^ 80'b00000000000000000000000000000010000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1011101100010100:begin data = code ^ 80'b00000000000000000000000000000010000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1101110001011110:begin data = code ^ 80'b00000000000000000000000000000010000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0001001011001010:begin data = code ^ 80'b00000000000000000000000000000010000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0000001000001111:begin data = code ^ 80'b00000000000000000000000000000010000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0010001110000101:begin data = code ^ 80'b00000000000000000000000000000010000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000010010001:begin data = code ^ 80'b00000000000000000000000000000010000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1110011010111001:begin data = code ^ 80'b00000000000000000000000000000010000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011100000100:begin data = code ^ 80'b00000000000000000000000000000010001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110100110010011:begin data = code ^ 80'b00000000000000000000000000000010010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111100101010000:begin data = code ^ 80'b00000000000000000000000000000010100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101010100111011:begin data = code ^ 80'b00000000000000000000000000000011000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111001001000:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1011111001001011:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1011111001001101:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1011111001000001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1011111001011001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1011111001101001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1011111000001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1011111011001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1011111101001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1011110001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1011101001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1011011001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1010111001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1001111001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1111111001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0011111001001001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0011001110100100:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0010100001111110:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0001111111001010:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0111000010100010:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1010111001110010:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1001111000111111:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1111111010100101:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0011111110010001:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0011000000010100:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0010111100011110:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0001000100001010:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0110110100100010:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1001010101110010:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1110100000111111:begin data = code ^ 80'b00000000000000000000000000000100000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0001001010100101:begin data = code ^ 80'b00000000000000000000000000000100000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0110101001111100:begin data = code ^ 80'b00000000000000000000000000000100000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1001101111001110:begin data = code ^ 80'b00000000000000000000000000000100000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1111010101000111:begin data = code ^ 80'b00000000000000000000000000000100000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0010100001010101:begin data = code ^ 80'b00000000000000000000000000000100000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0001111110011100:begin data = code ^ 80'b00000000000000000000000000000100000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0111000000001110:begin data = code ^ 80'b00000000000000000000000000000100000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1010111100101010:begin data = code ^ 80'b00000000000000000000000000000100000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1001110010001111:begin data = code ^ 80'b00000000000000000000000000000100000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1111101111000101:begin data = code ^ 80'b00000000000000000000000000000100000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0011010101010001:begin data = code ^ 80'b00000000000000000000000000000100000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0010010110010100:begin data = code ^ 80'b00000000000000000000000000000100000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0000010000011110:begin data = code ^ 80'b00000000000000000000000000000100000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011100001010:begin data = code ^ 80'b00000000000000000000000000000100000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1100000100100010:begin data = code ^ 80'b00000000000000000000000000000100000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0100000010011111:begin data = code ^ 80'b00000000000000000000000000000100001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111000001000:begin data = code ^ 80'b00000000000000000000000000000100010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111011001011:begin data = code ^ 80'b00000000000000000000000000000100100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111001010100000:begin data = code ^ 80'b00000000000000000000000000000101000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011110011011:begin data = code ^ 80'b00000000000000000000000000000110000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000101111110:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1111000101111101:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1111000101111011:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1111000101110111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1111000101101111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1111000101011111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1111000100111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1111000111111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1111000001111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1111001101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1111010101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1111100101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1110000101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1101000101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1011000101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0111000101111111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0111110010010010:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0110011101001000:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0101000011111100:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0011111110010100:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1110000101000100:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1101000100001001:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1011000110010011:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0111000010100111:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0111111100100010:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0110000000101000:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0101111000111100:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0010001000010100:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1101101001000100:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1010011100001001:begin data = code ^ 80'b00000000000000000000000000001000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0101110110010011:begin data = code ^ 80'b00000000000000000000000000001000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0010010101001010:begin data = code ^ 80'b00000000000000000000000000001000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1101010011111000:begin data = code ^ 80'b00000000000000000000000000001000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1011101001110001:begin data = code ^ 80'b00000000000000000000000000001000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0110011101100011:begin data = code ^ 80'b00000000000000000000000000001000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0101000010101010:begin data = code ^ 80'b00000000000000000000000000001000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0011111100111000:begin data = code ^ 80'b00000000000000000000000000001000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1110000000011100:begin data = code ^ 80'b00000000000000000000000000001000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1101001110111001:begin data = code ^ 80'b00000000000000000000000000001000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1011010011110011:begin data = code ^ 80'b00000000000000000000000000001000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0111101001100111:begin data = code ^ 80'b00000000000000000000000000001000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0110101010100010:begin data = code ^ 80'b00000000000000000000000000001000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0100101100101000:begin data = code ^ 80'b00000000000000000000000000001000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100000111100:begin data = code ^ 80'b00000000000000000000000000001000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111000010100:begin data = code ^ 80'b00000000000000000000000000001000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111110101001:begin data = code ^ 80'b00000000000000000000000000001000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000100111110:begin data = code ^ 80'b00000000000000000000000000001000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000111111101:begin data = code ^ 80'b00000000000000000000000000001000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110110010110:begin data = code ^ 80'b00000000000000000000000000001001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110100010101101:begin data = code ^ 80'b00000000000000000000000000001010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100111100110110:begin data = code ^ 80'b00000000000000000000000000001100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111100010010:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0110111100010001:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0110111100010111:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0110111100011011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0110111100000011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0110111100110011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0110111101010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0110111110010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0110111000010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0110110100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0110101100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0110011100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0111111100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0100111100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0010111100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1110111100010011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1110001011111110:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1111100100100100:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1100111010010000:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1010000111111000:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0111111100101000:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0100111101100101:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0010111111111111:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1110111011001011:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1110000101001110:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1111111001000100:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1100000001010000:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1011110001111000:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0100010000101000:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0011100101100101:begin data = code ^ 80'b00000000000000000000000000010000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1100001111111111:begin data = code ^ 80'b00000000000000000000000000010000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1011101100100110:begin data = code ^ 80'b00000000000000000000000000010000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0100101010010100:begin data = code ^ 80'b00000000000000000000000000010000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0010010000011101:begin data = code ^ 80'b00000000000000000000000000010000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1111100100001111:begin data = code ^ 80'b00000000000000000000000000010000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1100111011000110:begin data = code ^ 80'b00000000000000000000000000010000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1010000101010100:begin data = code ^ 80'b00000000000000000000000000010000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0111111001110000:begin data = code ^ 80'b00000000000000000000000000010000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0100110111010101:begin data = code ^ 80'b00000000000000000000000000010000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0010101010011111:begin data = code ^ 80'b00000000000000000000000000010000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1110010000001011:begin data = code ^ 80'b00000000000000000000000000010000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1111010011001110:begin data = code ^ 80'b00000000000000000000000000010000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1101010101000100:begin data = code ^ 80'b00000000000000000000000000010000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1001011001010000:begin data = code ^ 80'b00000000000000000000000000010000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000001111000:begin data = code ^ 80'b00000000000000000000000000010000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000111000101:begin data = code ^ 80'b00000000000000000000000000010000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001111101010010:begin data = code ^ 80'b00000000000000000000000000010000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111110010001:begin data = code ^ 80'b00000000000000000000000000010000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010001111111010:begin data = code ^ 80'b00000000000000000000000000010001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011011000001:begin data = code ^ 80'b00000000000000000000000000010010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000101011010:begin data = code ^ 80'b00000000000000000000000000010100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001111001101100:begin data = code ^ 80'b00000000000000000000000000011000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111000100111:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1101111000100100:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1101111000100010:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1101111000101110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1101111000110110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1101111000000110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1101111001100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1101111010100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1101111100100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1101110000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1101101000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1101011000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1100111000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1111111000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1001111000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0101111000100110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0101001111001011:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0100100000010001:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0111111110100101:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0001000011001101:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1100111000011101:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1111111001010000:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1001111011001010:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0101111111111110:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0101000001111011:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0100111101110001:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0111000101100101:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0000110101001101:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1111010100011101:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1000100001010000:begin data = code ^ 80'b00000000000000000000000000100000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0111001011001010:begin data = code ^ 80'b00000000000000000000000000100000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0000101000010011:begin data = code ^ 80'b00000000000000000000000000100000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1111101110100001:begin data = code ^ 80'b00000000000000000000000000100000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1001010100101000:begin data = code ^ 80'b00000000000000000000000000100000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0100100000111010:begin data = code ^ 80'b00000000000000000000000000100000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0111111111110011:begin data = code ^ 80'b00000000000000000000000000100000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0001000001100001:begin data = code ^ 80'b00000000000000000000000000100000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1100111101000101:begin data = code ^ 80'b00000000000000000000000000100000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1111110011100000:begin data = code ^ 80'b00000000000000000000000000100000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1001101110101010:begin data = code ^ 80'b00000000000000000000000000100000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0101010100111110:begin data = code ^ 80'b00000000000000000000000000100000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0100010111111011:begin data = code ^ 80'b00000000000000000000000000100000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0110010001110001:begin data = code ^ 80'b00000000000000000000000000100000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011101100101:begin data = code ^ 80'b00000000000000000000000000100000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000101001101:begin data = code ^ 80'b00000000000000000000000000100000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000011110000:begin data = code ^ 80'b00000000000000000000000000100000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111001100111:begin data = code ^ 80'b00000000000000000000000000100000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111010100100:begin data = code ^ 80'b00000000000000000000000000100000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001011001111:begin data = code ^ 80'b00000000000000000000000000100001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011111110100:begin data = code ^ 80'b00000000000000000000000000100010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000001101111:begin data = code ^ 80'b00000000000000000000000000100100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111101011001:begin data = code ^ 80'b00000000000000000000000000101000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011000100110101:begin data = code ^ 80'b00000000000000000000000000110000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000110100000:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0011000110100011:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0011000110100101:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0011000110101001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0011000110110001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0011000110000001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0011000111100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0011000100100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0011000010100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0011001110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0011010110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0011100110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0010000110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0001000110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0111000110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1011000110100001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1011110001001100:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1010011110010110:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1001000000100010:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1111111101001010:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0010000110011010:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0001000111010111:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0111000101001101:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1011000001111001:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1011111111111100:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1010000011110110:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1001111011100010:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1110001011001010:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0001101010011010:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0110011111010111:begin data = code ^ 80'b00000000000000000000000001000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1001110101001101:begin data = code ^ 80'b00000000000000000000000001000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1110010110010100:begin data = code ^ 80'b00000000000000000000000001000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0001010000100110:begin data = code ^ 80'b00000000000000000000000001000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0111101010101111:begin data = code ^ 80'b00000000000000000000000001000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1010011110111101:begin data = code ^ 80'b00000000000000000000000001000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1001000001110100:begin data = code ^ 80'b00000000000000000000000001000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1111111111100110:begin data = code ^ 80'b00000000000000000000000001000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0010000011000010:begin data = code ^ 80'b00000000000000000000000001000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0001001101100111:begin data = code ^ 80'b00000000000000000000000001000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0111010000101101:begin data = code ^ 80'b00000000000000000000000001000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1011101010111001:begin data = code ^ 80'b00000000000000000000000001000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1010101001111100:begin data = code ^ 80'b00000000000000000000000001000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1000101111110110:begin data = code ^ 80'b00000000000000000000000001000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100011100010:begin data = code ^ 80'b00000000000000000000000001000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0100111011001010:begin data = code ^ 80'b00000000000000000000000001000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111101110111:begin data = code ^ 80'b00000000000000000000000001000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100000111100000:begin data = code ^ 80'b00000000000000000000000001000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000100100011:begin data = code ^ 80'b00000000000000000000000001000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111110101001000:begin data = code ^ 80'b00000000000000000000000001000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100001110011:begin data = code ^ 80'b00000000000000000000000001000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111111101000:begin data = code ^ 80'b00000000000000000000000001000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100000011011110:begin data = code ^ 80'b00000000000000000000000001001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111010110010:begin data = code ^ 80'b00000000000000000000000001010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111110000111:begin data = code ^ 80'b00000000000000000000000001100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001101000011:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0110001101000000:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0110001101000110:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0110001101001010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0110001101010010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0110001101100010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0110001100000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0110001111000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0110001001000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0110000101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0110011101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0110101101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0111001101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0100001101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0010001101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1110001101000010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1110111010101111:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1111010101110101:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1100001011000001:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1010110110101001:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0111001101111001:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0100001100110100:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0010001110101110:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1110001010011010:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1110110100011111:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1111001000010101:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1100110000000001:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1011000000101001:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0100100001111001:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0011010100110100:begin data = code ^ 80'b00000000000000000000000010000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1100111110101110:begin data = code ^ 80'b00000000000000000000000010000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1011011101110111:begin data = code ^ 80'b00000000000000000000000010000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0100011011000101:begin data = code ^ 80'b00000000000000000000000010000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0010100001001100:begin data = code ^ 80'b00000000000000000000000010000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1111010101011110:begin data = code ^ 80'b00000000000000000000000010000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1100001010010111:begin data = code ^ 80'b00000000000000000000000010000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1010110100000101:begin data = code ^ 80'b00000000000000000000000010000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0111001000100001:begin data = code ^ 80'b00000000000000000000000010000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0100000110000100:begin data = code ^ 80'b00000000000000000000000010000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0010011011001110:begin data = code ^ 80'b00000000000000000000000010000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1110100001011010:begin data = code ^ 80'b00000000000000000000000010000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1111100010011111:begin data = code ^ 80'b00000000000000000000000010000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1101100100010101:begin data = code ^ 80'b00000000000000000000000010000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1001101000000001:begin data = code ^ 80'b00000000000000000000000010000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110000101001:begin data = code ^ 80'b00000000000000000000000010000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1001110110010100:begin data = code ^ 80'b00000000000000000000000010000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001100000011:begin data = code ^ 80'b00000000000000000000000010000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000001111000000:begin data = code ^ 80'b00000000000000000000000010000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111110101011:begin data = code ^ 80'b00000000000000000000000010000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111101010010000:begin data = code ^ 80'b00000000000000000000000010000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101110100001011:begin data = code ^ 80'b00000000000000000000000010000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001000111101:begin data = code ^ 80'b00000000000000000000000010001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000110001010001:begin data = code ^ 80'b00000000000000000000000010010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110101100100:begin data = code ^ 80'b00000000000000000000000010100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101001011100011:begin data = code ^ 80'b00000000000000000000000011000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011010000101:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1100011010000110:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1100011010000000:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1100011010001100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1100011010010100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1100011010100100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1100011011000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1100011000000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1100011110000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1100010010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1100001010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1100111010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1101011010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1110011010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1000011010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0100011010000100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0100101101101001:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0101000010110011:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0110011100000111:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0000100001101111:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1101011010111111:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1110011011110010:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1000011001101000:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0100011101011100:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0100100011011001:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0101011111010011:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0110100111000111:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0001010111101111:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1110110110111111:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1001000011110010:begin data = code ^ 80'b00000000000000000000000100000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0110101001101000:begin data = code ^ 80'b00000000000000000000000100000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0001001010110001:begin data = code ^ 80'b00000000000000000000000100000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1110001100000011:begin data = code ^ 80'b00000000000000000000000100000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1000110110001010:begin data = code ^ 80'b00000000000000000000000100000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0101000010011000:begin data = code ^ 80'b00000000000000000000000100000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0110011101010001:begin data = code ^ 80'b00000000000000000000000100000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0000100011000011:begin data = code ^ 80'b00000000000000000000000100000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1101011111100111:begin data = code ^ 80'b00000000000000000000000100000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1110010001000010:begin data = code ^ 80'b00000000000000000000000100000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1000001100001000:begin data = code ^ 80'b00000000000000000000000100000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0100110110011100:begin data = code ^ 80'b00000000000000000000000100000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0101110101011001:begin data = code ^ 80'b00000000000000000000000100000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0111110011010011:begin data = code ^ 80'b00000000000000000000000100000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111111000111:begin data = code ^ 80'b00000000000000000000000100000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1011100111101111:begin data = code ^ 80'b00000000000000000000000100000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100001010010:begin data = code ^ 80'b00000000000000000000000100000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011011011000101:begin data = code ^ 80'b00000000000000000000000100000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011000000110:begin data = code ^ 80'b00000000000000000000000100000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101001101101:begin data = code ^ 80'b00000000000000000000000100000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111101010110:begin data = code ^ 80'b00000000000000000000000100000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111100011001101:begin data = code ^ 80'b00000000000000000000000100000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011011111111011:begin data = code ^ 80'b00000000000000000000000100001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100110010111:begin data = code ^ 80'b00000000000000000000000100010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100010100010:begin data = code ^ 80'b00000000000000000000000100100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011100100101:begin data = code ^ 80'b00000000000000000000000101000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010010111000110:begin data = code ^ 80'b00000000000000000000000110000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000011100100:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0000000011100111:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0000000011100001:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0000000011101101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0000000011110101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0000000011000101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0000000010100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0000000001100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0000000111100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0000001011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0000010011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0000100011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0001000011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0010000011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0100000011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1000000011100101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1000110100001000:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1001011011010010:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1010000101100110:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1100111000001110:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0001000011011110:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0010000010010011:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0100000000001001:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1000000100111101:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1000111010111000:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1001000110110010:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1010111110100110:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1101001110001110:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0010101111011110:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0101011010010011:begin data = code ^ 80'b00000000000000000000001000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1010110000001001:begin data = code ^ 80'b00000000000000000000001000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1101010011010000:begin data = code ^ 80'b00000000000000000000001000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0010010101100010:begin data = code ^ 80'b00000000000000000000001000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0100101111101011:begin data = code ^ 80'b00000000000000000000001000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1001011011111001:begin data = code ^ 80'b00000000000000000000001000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1010000100110000:begin data = code ^ 80'b00000000000000000000001000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1100111010100010:begin data = code ^ 80'b00000000000000000000001000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0001000110000110:begin data = code ^ 80'b00000000000000000000001000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0010001000100011:begin data = code ^ 80'b00000000000000000000001000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0100010101101001:begin data = code ^ 80'b00000000000000000000001000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1000101111111101:begin data = code ^ 80'b00000000000000000000001000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1001101100111000:begin data = code ^ 80'b00000000000000000000001000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1011101010110010:begin data = code ^ 80'b00000000000000000000001000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100110100110:begin data = code ^ 80'b00000000000000000000001000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111110001110:begin data = code ^ 80'b00000000000000000000001000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111000110011:begin data = code ^ 80'b00000000000000000000001000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000010100100:begin data = code ^ 80'b00000000000000000000001000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000001100111:begin data = code ^ 80'b00000000000000000000001000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110000001100:begin data = code ^ 80'b00000000000000000000001000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100100110111:begin data = code ^ 80'b00000000000000000000001000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111010101100:begin data = code ^ 80'b00000000000000000000001000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000110011010:begin data = code ^ 80'b00000000000000000000001000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111111110110:begin data = code ^ 80'b00000000000000000000001000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111011000011:begin data = code ^ 80'b00000000000000000000001000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000101000100:begin data = code ^ 80'b00000000000000000000001001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001110100111:begin data = code ^ 80'b00000000000000000000001010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011001100001:begin data = code ^ 80'b00000000000000000000001100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000111001011:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0000000111001000:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0000000111001110:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0000000111000010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0000000111011010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0000000111101010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0000000110001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0000000101001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0000000011001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0000001111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0000010111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0000100111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0001000111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0010000111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0100000111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1000000111001010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1000110000100111:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1001011111111101:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1010000001001001:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1100111100100001:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0001000111110001:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0010000110111100:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0100000100100110:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1000000000010010:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1000111110010111:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1001000010011101:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1010111010001001:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1101001010100001:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0010101011110001:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0101011110111100:begin data = code ^ 80'b00000000000000000000010000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1010110100100110:begin data = code ^ 80'b00000000000000000000010000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1101010111111111:begin data = code ^ 80'b00000000000000000000010000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0010010001001101:begin data = code ^ 80'b00000000000000000000010000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0100101011000100:begin data = code ^ 80'b00000000000000000000010000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1001011111010110:begin data = code ^ 80'b00000000000000000000010000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1010000000011111:begin data = code ^ 80'b00000000000000000000010000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1100111110001101:begin data = code ^ 80'b00000000000000000000010000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0001000010101001:begin data = code ^ 80'b00000000000000000000010000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0010001100001100:begin data = code ^ 80'b00000000000000000000010000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0100010001000110:begin data = code ^ 80'b00000000000000000000010000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1000101011010010:begin data = code ^ 80'b00000000000000000000010000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1001101000010111:begin data = code ^ 80'b00000000000000000000010000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1011101110011101:begin data = code ^ 80'b00000000000000000000010000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100010001001:begin data = code ^ 80'b00000000000000000000010000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111010100001:begin data = code ^ 80'b00000000000000000000010000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111100011100:begin data = code ^ 80'b00000000000000000000010000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000110001011:begin data = code ^ 80'b00000000000000000000010000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000101001000:begin data = code ^ 80'b00000000000000000000010000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110100100011:begin data = code ^ 80'b00000000000000000000010000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100000011000:begin data = code ^ 80'b00000000000000000000010000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111110000011:begin data = code ^ 80'b00000000000000000000010000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000010110101:begin data = code ^ 80'b00000000000000000000010000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111011011001:begin data = code ^ 80'b00000000000000000000010000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111111101100:begin data = code ^ 80'b00000000000000000000010000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000001101011:begin data = code ^ 80'b00000000000000000000010001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001010001000:begin data = code ^ 80'b00000000000000000000010010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011101001110:begin data = code ^ 80'b00000000000000000000010100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000100101111:begin data = code ^ 80'b00000000000000000000011000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001110010101:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0000001110010110:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0000001110010000:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0000001110011100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0000001110000100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0000001110110100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0000001111010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0000001100010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0000001010010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0000000110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0000011110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0000101110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0001001110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0010001110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0100001110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1000001110010100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1000111001111001:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1001010110100011:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1010001000010111:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1100110101111111:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0001001110101111:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0010001111100010:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0100001101111000:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1000001001001100:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1000110111001001:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1001001011000011:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1010110011010111:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1101000011111111:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0010100010101111:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0101010111100010:begin data = code ^ 80'b00000000000000000000100000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1010111101111000:begin data = code ^ 80'b00000000000000000000100000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1101011110100001:begin data = code ^ 80'b00000000000000000000100000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0010011000010011:begin data = code ^ 80'b00000000000000000000100000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0100100010011010:begin data = code ^ 80'b00000000000000000000100000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1001010110001000:begin data = code ^ 80'b00000000000000000000100000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1010001001000001:begin data = code ^ 80'b00000000000000000000100000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1100110111010011:begin data = code ^ 80'b00000000000000000000100000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0001001011110111:begin data = code ^ 80'b00000000000000000000100000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0010000101010010:begin data = code ^ 80'b00000000000000000000100000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0100011000011000:begin data = code ^ 80'b00000000000000000000100000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1000100010001100:begin data = code ^ 80'b00000000000000000000100000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1001100001001001:begin data = code ^ 80'b00000000000000000000100000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1011100111000011:begin data = code ^ 80'b00000000000000000000100000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1111101011010111:begin data = code ^ 80'b00000000000000000000100000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0111110011111111:begin data = code ^ 80'b00000000000000000000100000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1111110101000010:begin data = code ^ 80'b00000000000000000000100000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001111010101:begin data = code ^ 80'b00000000000000000000100000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001100010110:begin data = code ^ 80'b00000000000000000000100000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100111101111101:begin data = code ^ 80'b00000000000000000000100000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001101001000110:begin data = code ^ 80'b00000000000000000000100000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110111011101:begin data = code ^ 80'b00000000000000000000100000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111001011101011:begin data = code ^ 80'b00000000000000000000100000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110110010000111:begin data = code ^ 80'b00000000000000000000100000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101110110110010:begin data = code ^ 80'b00000000000000000000100000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001000110101:begin data = code ^ 80'b00000000000000000000100001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000011010110:begin data = code ^ 80'b00000000000000000000100010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100010100010000:begin data = code ^ 80'b00000000000000000000100100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001101110001:begin data = code ^ 80'b00000000000000000000101000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001001011110:begin data = code ^ 80'b00000000000000000000110000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011100101001:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0000011100101010:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0000011100101100:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0000011100100000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0000011100111000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0000011100001000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0000011101101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0000011110101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0000011000101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0000010100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0000001100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0000111100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0001011100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0010011100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0100011100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1000011100101000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1000101011000101:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1001000100011111:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1010011010101011:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1100100111000011:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0001011100010011:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0010011101011110:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0100011111000100:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1000011011110000:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1000100101110101:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1001011001111111:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1010100001101011:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1101010001000011:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0010110000010011:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0101000101011110:begin data = code ^ 80'b00000000000000000001000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1010101111000100:begin data = code ^ 80'b00000000000000000001000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1101001100011101:begin data = code ^ 80'b00000000000000000001000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0010001010101111:begin data = code ^ 80'b00000000000000000001000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0100110000100110:begin data = code ^ 80'b00000000000000000001000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1001000100110100:begin data = code ^ 80'b00000000000000000001000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1010011011111101:begin data = code ^ 80'b00000000000000000001000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1100100101101111:begin data = code ^ 80'b00000000000000000001000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0001011001001011:begin data = code ^ 80'b00000000000000000001000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0010010111101110:begin data = code ^ 80'b00000000000000000001000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0100001010100100:begin data = code ^ 80'b00000000000000000001000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1000110000110000:begin data = code ^ 80'b00000000000000000001000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1001110011110101:begin data = code ^ 80'b00000000000000000001000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1011110101111111:begin data = code ^ 80'b00000000000000000001000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111001101011:begin data = code ^ 80'b00000000000000000001000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0111100001000011:begin data = code ^ 80'b00000000000000000001000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100111111110:begin data = code ^ 80'b00000000000000000001000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011101101001:begin data = code ^ 80'b00000000000000000001000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110011110101010:begin data = code ^ 80'b00000000000000000001000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100101111000001:begin data = code ^ 80'b00000000000000000001000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001111011111010:begin data = code ^ 80'b00000000000000000001000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011100101100001:begin data = code ^ 80'b00000000000000000001000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011001010111:begin data = code ^ 80'b00000000000000000001000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110100000111011:begin data = code ^ 80'b00000000000000000001000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101100100001110:begin data = code ^ 80'b00000000000000000001000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011011010001001:begin data = code ^ 80'b00000000000000000001000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110010001101010:begin data = code ^ 80'b00000000000000000001000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100000110101100:begin data = code ^ 80'b00000000000000000001000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011111001101:begin data = code ^ 80'b00000000000000000001001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011011100010:begin data = code ^ 80'b00000000000000000001010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000010010111100:begin data = code ^ 80'b00000000000000000001100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111001010001:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0000111001010010:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0000111001010100:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0000111001011000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0000111001000000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0000111001110000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0000111000010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0000111011010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0000111101010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0000110001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0000101001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0000011001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0001111001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0010111001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0100111001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1000111001010000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1000001110111101:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1001100001100111:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1010111111010011:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1100000010111011:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0001111001101011:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0010111000100110:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0100111010111100:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1000111110001000:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1000000000001101:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1001111100000111:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1010000100010011:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1101110100111011:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0010010101101011:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0101100000100110:begin data = code ^ 80'b00000000000000000010000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1010001010111100:begin data = code ^ 80'b00000000000000000010000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1101101001100101:begin data = code ^ 80'b00000000000000000010000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0010101111010111:begin data = code ^ 80'b00000000000000000010000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0100010101011110:begin data = code ^ 80'b00000000000000000010000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1001100001001100:begin data = code ^ 80'b00000000000000000010000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1010111110000101:begin data = code ^ 80'b00000000000000000010000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1100000000010111:begin data = code ^ 80'b00000000000000000010000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0001111100110011:begin data = code ^ 80'b00000000000000000010000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0010110010010110:begin data = code ^ 80'b00000000000000000010000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0100101111011100:begin data = code ^ 80'b00000000000000000010000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1000010101001000:begin data = code ^ 80'b00000000000000000010000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1001010110001101:begin data = code ^ 80'b00000000000000000010000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1011010000000111:begin data = code ^ 80'b00000000000000000010000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011100010011:begin data = code ^ 80'b00000000000000000010000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000100111011:begin data = code ^ 80'b00000000000000000010000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000010000110:begin data = code ^ 80'b00000000000000000010000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111000010001:begin data = code ^ 80'b00000000000000000010000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111011010010:begin data = code ^ 80'b00000000000000000010000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001010111001:begin data = code ^ 80'b00000000000000000010000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001011110000010:begin data = code ^ 80'b00000000000000000010000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011000000011001:begin data = code ^ 80'b00000000000000000010000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111100101111:begin data = code ^ 80'b00000000000000000010000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000101000011:begin data = code ^ 80'b00000000000000000010000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000001110110:begin data = code ^ 80'b00000000000000000010000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111111110001:begin data = code ^ 80'b00000000000000000010000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110110100010010:begin data = code ^ 80'b00000000000000000010000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100011010100:begin data = code ^ 80'b00000000000000000010000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111010110101:begin data = code ^ 80'b00000000000000000010001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111110011010:begin data = code ^ 80'b00000000000000000010010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000110111000100:begin data = code ^ 80'b00000000000000000010100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100101111000:begin data = code ^ 80'b00000000000000000011000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110010100001:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0001110010100010:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0001110010100100:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0001110010101000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0001110010110000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0001110010000000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0001110011100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0001110000100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0001110110100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0001111010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0001100010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0001010010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0000110010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0011110010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0101110010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1001110010100000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1001000101001101:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1000101010010111:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1011110100100011:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1101001001001011:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0000110010011011:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0011110011010110:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0101110001001100:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1001110101111000:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1001001011111101:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1000110111110111:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1011001111100011:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1100111111001011:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0011011110011011:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0100101011010110:begin data = code ^ 80'b00000000000000000100000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1011000001001100:begin data = code ^ 80'b00000000000000000100000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1100100010010101:begin data = code ^ 80'b00000000000000000100000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0011100100100111:begin data = code ^ 80'b00000000000000000100000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0101011110101110:begin data = code ^ 80'b00000000000000000100000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1000101010111100:begin data = code ^ 80'b00000000000000000100000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1011110101110101:begin data = code ^ 80'b00000000000000000100000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1101001011100111:begin data = code ^ 80'b00000000000000000100000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0000110111000011:begin data = code ^ 80'b00000000000000000100000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0011111001100110:begin data = code ^ 80'b00000000000000000100000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0101100100101100:begin data = code ^ 80'b00000000000000000100000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1001011110111000:begin data = code ^ 80'b00000000000000000100000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1000011101111101:begin data = code ^ 80'b00000000000000000100000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1010011011110111:begin data = code ^ 80'b00000000000000000100000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010111100011:begin data = code ^ 80'b00000000000000000100000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001111001011:begin data = code ^ 80'b00000000000000000100000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001001110110:begin data = code ^ 80'b00000000000000000100000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110110011100001:begin data = code ^ 80'b00000000000000000100000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111110000100010:begin data = code ^ 80'b00000000000000000100000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000001001001:begin data = code ^ 80'b00000000000000000100000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010101110010:begin data = code ^ 80'b00000000000000000100000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010001011101001:begin data = code ^ 80'b00000000000000000100000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110110111011111:begin data = code ^ 80'b00000000000000000100000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001110110011:begin data = code ^ 80'b00000000000000000100000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001010000110:begin data = code ^ 80'b00000000000000000100000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110100000001:begin data = code ^ 80'b00000000000000000100000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111111100010:begin data = code ^ 80'b00000000000000000100000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101101000100100:begin data = code ^ 80'b00000000000000000100000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110001000101:begin data = code ^ 80'b00000000000000000100001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110101101010:begin data = code ^ 80'b00000000000000000100010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001111100110100:begin data = code ^ 80'b00000000000000000100100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001101110001000:begin data = code ^ 80'b00000000000000000101000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001011110000:begin data = code ^ 80'b00000000000000000110000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100101000001:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0011100101000010:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0011100101000100:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0011100101001000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0011100101010000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0011100101100000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0011100100000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0011100111000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0011100001000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0011101101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0011110101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0011000101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0010100101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0001100101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0111100101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1011100101000000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1011010010101101:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1010111101110111:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1001100011000011:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1111011110101011:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0010100101111011:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0001100100110110:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0111100110101100:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1011100010011000:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1011011100011101:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1010100000010111:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1001011000000011:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1110101000101011:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0001001001111011:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0110111100110110:begin data = code ^ 80'b00000000000000001000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1001010110101100:begin data = code ^ 80'b00000000000000001000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1110110101110101:begin data = code ^ 80'b00000000000000001000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0001110011000111:begin data = code ^ 80'b00000000000000001000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0111001001001110:begin data = code ^ 80'b00000000000000001000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1010111101011100:begin data = code ^ 80'b00000000000000001000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1001100010010101:begin data = code ^ 80'b00000000000000001000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1111011100000111:begin data = code ^ 80'b00000000000000001000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0010100000100011:begin data = code ^ 80'b00000000000000001000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0001101110000110:begin data = code ^ 80'b00000000000000001000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0111110011001100:begin data = code ^ 80'b00000000000000001000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1011001001011000:begin data = code ^ 80'b00000000000000001000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1010001010011101:begin data = code ^ 80'b00000000000000001000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1000001100010111:begin data = code ^ 80'b00000000000000001000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1100000000000011:begin data = code ^ 80'b00000000000000001000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011000101011:begin data = code ^ 80'b00000000000000001000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011110010110:begin data = code ^ 80'b00000000000000001000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100100000001:begin data = code ^ 80'b00000000000000001000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101100111000010:begin data = code ^ 80'b00000000000000001000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111010110101001:begin data = code ^ 80'b00000000000000001000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000010010010:begin data = code ^ 80'b00000000000000001000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011100001001:begin data = code ^ 80'b00000000000000001000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100000111111:begin data = code ^ 80'b00000000000000001000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101011001010011:begin data = code ^ 80'b00000000000000001000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110011101100110:begin data = code ^ 80'b00000000000000001000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100011100001:begin data = code ^ 80'b00000000000000001000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101101000000010:begin data = code ^ 80'b00000000000000001000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111111000100:begin data = code ^ 80'b00000000000000001000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100110100101:begin data = code ^ 80'b00000000000000001000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100010001010:begin data = code ^ 80'b00000000000000001000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011101011010100:begin data = code ^ 80'b00000000000000001000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111001101000:begin data = code ^ 80'b00000000000000001001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011011100010000:begin data = code ^ 80'b00000000000000001010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010010111100000:begin data = code ^ 80'b00000000000000001100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001010000001:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0111001010000010:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0111001010000100:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0111001010001000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0111001010010000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0111001010100000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0111001011000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0111001000000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0111001110000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0111000010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0111011010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0111101010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0110001010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0101001010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0011001010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1111001010000000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1111111101101101:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1110010010110111:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1101001100000011:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1011110001101011:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0110001010111011:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0101001011110110:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0011001001101100:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1111001101011000:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1111110011011101:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1110001111010111:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1101110111000011:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1010000111101011:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0101100110111011:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0010010011110110:begin data = code ^ 80'b00000000000000010000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1101111001101100:begin data = code ^ 80'b00000000000000010000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1010011010110101:begin data = code ^ 80'b00000000000000010000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0101011100000111:begin data = code ^ 80'b00000000000000010000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0011100110001110:begin data = code ^ 80'b00000000000000010000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1110010010011100:begin data = code ^ 80'b00000000000000010000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1101001101010101:begin data = code ^ 80'b00000000000000010000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1011110011000111:begin data = code ^ 80'b00000000000000010000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0110001111100011:begin data = code ^ 80'b00000000000000010000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0101000001000110:begin data = code ^ 80'b00000000000000010000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0011011100001100:begin data = code ^ 80'b00000000000000010000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1111100110011000:begin data = code ^ 80'b00000000000000010000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1110100101011101:begin data = code ^ 80'b00000000000000010000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1100100011010111:begin data = code ^ 80'b00000000000000010000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101111000011:begin data = code ^ 80'b00000000000000010000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0000110111101011:begin data = code ^ 80'b00000000000000010000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1000110001010110:begin data = code ^ 80'b00000000000000010000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001011000001:begin data = code ^ 80'b00000000000000010000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001000000010:begin data = code ^ 80'b00000000000000010000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111001101001:begin data = code ^ 80'b00000000000000010000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110101101010010:begin data = code ^ 80'b00000000000000010000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110011001001:begin data = code ^ 80'b00000000000000010000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000001111111111:begin data = code ^ 80'b00000000000000010000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110110010011:begin data = code ^ 80'b00000000000000010000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010110010100110:begin data = code ^ 80'b00000000000000010000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001100100001:begin data = code ^ 80'b00000000000000010000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000111000010:begin data = code ^ 80'b00000000000000010000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011010000000100:begin data = code ^ 80'b00000000000000010000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001001100101:begin data = code ^ 80'b00000000000000010000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001101001010:begin data = code ^ 80'b00000000000000010000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000100010100:begin data = code ^ 80'b00000000000000010000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111010110101000:begin data = code ^ 80'b00000000000000010001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111110011010000:begin data = code ^ 80'b00000000000000010010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111000100000:begin data = code ^ 80'b00000000000000010100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100101111000000:begin data = code ^ 80'b00000000000000011000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010100000001:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1110010100000010:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1110010100000100:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1110010100001000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1110010100010000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1110010100100000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1110010101000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1110010110000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1110010000000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1110011100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1110000100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1110110100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1111010100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1100010100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1010010100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0110010100000000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0110100011101101:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0111001100110111:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0100010010000011:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0010101111101011:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1111010100111011:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1100010101110110:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1010010111101100:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0110010011011000:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0110101101011101:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0111010001010111:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0100101001000011:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0011011001101011:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1100111000111011:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1011001101110110:begin data = code ^ 80'b00000000000000100000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0100100111101100:begin data = code ^ 80'b00000000000000100000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0011000100110101:begin data = code ^ 80'b00000000000000100000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1100000010000111:begin data = code ^ 80'b00000000000000100000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1010111000001110:begin data = code ^ 80'b00000000000000100000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0111001100011100:begin data = code ^ 80'b00000000000000100000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0100010011010101:begin data = code ^ 80'b00000000000000100000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0010101101000111:begin data = code ^ 80'b00000000000000100000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1111010001100011:begin data = code ^ 80'b00000000000000100000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1100011111000110:begin data = code ^ 80'b00000000000000100000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1010000010001100:begin data = code ^ 80'b00000000000000100000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0110111000011000:begin data = code ^ 80'b00000000000000100000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0111111011011101:begin data = code ^ 80'b00000000000000100000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0101111101010111:begin data = code ^ 80'b00000000000000100000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110001000011:begin data = code ^ 80'b00000000000000100000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1001101001101011:begin data = code ^ 80'b00000000000000100000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0001101111010110:begin data = code ^ 80'b00000000000000100000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001010101000001:begin data = code ^ 80'b00000000000000100000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000010110000010:begin data = code ^ 80'b00000000000000100000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100111101001:begin data = code ^ 80'b00000000000000100000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111110011010010:begin data = code ^ 80'b00000000000000100000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101101101001001:begin data = code ^ 80'b00000000000000100000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001010001111111:begin data = code ^ 80'b00000000000000100000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101000010011:begin data = code ^ 80'b00000000000000100000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011101100100110:begin data = code ^ 80'b00000000000000100000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101010010100001:begin data = code ^ 80'b00000000000000100000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011001000010:begin data = code ^ 80'b00000000000000100000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010001110000100:begin data = code ^ 80'b00000000000000100000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010111100101:begin data = code ^ 80'b00000000000000100000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010011001010:begin data = code ^ 80'b00000000000000100000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110011010010100:begin data = code ^ 80'b00000000000000100000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001000101000:begin data = code ^ 80'b00000000000000100001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110101101010000:begin data = code ^ 80'b00000000000000100010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100110100000:begin data = code ^ 80'b00000000000000100100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101110001000000:begin data = code ^ 80'b00000000000000101000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001011110000000:begin data = code ^ 80'b00000000000000110000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011111101100:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0100011111101111:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0100011111101001:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0100011111100101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0100011111111101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0100011111001101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0100011110101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0100011101101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0100011011101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0100010111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0100001111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0100111111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0101011111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0110011111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0000011111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1100011111101101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1100101000000000:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1101000111011010:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1110011001101110:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1000100100000110:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0101011111010110:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0110011110011011:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0000011100000001:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1100011000110101:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1100100110110000:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1101011010111010:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1110100010101110:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1001010010000110:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0110110011010110:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0001000110011011:begin data = code ^ 80'b00000000000001000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1110101100000001:begin data = code ^ 80'b00000000000001000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1001001111011000:begin data = code ^ 80'b00000000000001000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0110001001101010:begin data = code ^ 80'b00000000000001000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0000110011100011:begin data = code ^ 80'b00000000000001000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1101000111110001:begin data = code ^ 80'b00000000000001000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1110011000111000:begin data = code ^ 80'b00000000000001000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1000100110101010:begin data = code ^ 80'b00000000000001000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0101011010001110:begin data = code ^ 80'b00000000000001000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0110010100101011:begin data = code ^ 80'b00000000000001000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0000001001100001:begin data = code ^ 80'b00000000000001000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1100110011110101:begin data = code ^ 80'b00000000000001000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1101110000110000:begin data = code ^ 80'b00000000000001000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1111110110111010:begin data = code ^ 80'b00000000000001000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111010101110:begin data = code ^ 80'b00000000000001000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100010000110:begin data = code ^ 80'b00000000000001000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1011100100111011:begin data = code ^ 80'b00000000000001000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011011110101100:begin data = code ^ 80'b00000000000001000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010011101101111:begin data = code ^ 80'b00000000000001000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101100000100:begin data = code ^ 80'b00000000000001000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111000111111:begin data = code ^ 80'b00000000000001000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100110100100:begin data = code ^ 80'b00000000000001000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011011010010010:begin data = code ^ 80'b00000000000001000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010100011111110:begin data = code ^ 80'b00000000000001000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100111001011:begin data = code ^ 80'b00000000000001000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011001001100:begin data = code ^ 80'b00000000000001000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010010010101111:begin data = code ^ 80'b00000000000001000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000101101001:begin data = code ^ 80'b00000000000001000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011100001000:begin data = code ^ 80'b00000000000001000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011000100111:begin data = code ^ 80'b00000000000001000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100010001111001:begin data = code ^ 80'b00000000000001000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100000011000101:begin data = code ^ 80'b00000000000001000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100110111101:begin data = code ^ 80'b00000000000001000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101101101001101:begin data = code ^ 80'b00000000000001000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111010101101:begin data = code ^ 80'b00000000000001001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011010101101101:begin data = code ^ 80'b00000000000001010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010001011101101:begin data = code ^ 80'b00000000000001100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111111011011:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1000111111011000:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1000111111011110:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1000111111010010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1000111111001010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1000111111111010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1000111110011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1000111101011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1000111011011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1000110111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1000101111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1000011111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1001111111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1010111111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1100111111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0000111111011010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0000001000110111:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0001100111101101:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0010111001011001:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0100000100110001:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1001111111100001:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1010111110101100:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1100111100110110:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0000111000000010:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0000000110000111:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0001111010001101:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0010000010011001:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0101110010110001:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1010010011100001:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1101100110101100:begin data = code ^ 80'b00000000000010000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0010001100110110:begin data = code ^ 80'b00000000000010000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0101101111101111:begin data = code ^ 80'b00000000000010000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1010101001011101:begin data = code ^ 80'b00000000000010000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1100010011010100:begin data = code ^ 80'b00000000000010000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0001100111000110:begin data = code ^ 80'b00000000000010000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0010111000001111:begin data = code ^ 80'b00000000000010000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0100000110011101:begin data = code ^ 80'b00000000000010000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1001111010111001:begin data = code ^ 80'b00000000000010000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1010110100011100:begin data = code ^ 80'b00000000000010000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1100101001010110:begin data = code ^ 80'b00000000000010000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0000010011000010:begin data = code ^ 80'b00000000000010000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0001010000000111:begin data = code ^ 80'b00000000000010000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0011010110001101:begin data = code ^ 80'b00000000000010000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011010011001:begin data = code ^ 80'b00000000000010000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000010110001:begin data = code ^ 80'b00000000000010000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000100001100:begin data = code ^ 80'b00000000000010000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111110011011:begin data = code ^ 80'b00000000000010000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111101011000:begin data = code ^ 80'b00000000000010000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001100110011:begin data = code ^ 80'b00000000000010000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011000001000:begin data = code ^ 80'b00000000000010000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000110010011:begin data = code ^ 80'b00000000000010000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111010100101:begin data = code ^ 80'b00000000000010000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000011001001:begin data = code ^ 80'b00000000000010000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000111111100:begin data = code ^ 80'b00000000000010000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111001111011:begin data = code ^ 80'b00000000000010000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110110010011000:begin data = code ^ 80'b00000000000010000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100101011110:begin data = code ^ 80'b00000000000010000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111100111111:begin data = code ^ 80'b00000000000010000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111000010000:begin data = code ^ 80'b00000000000010000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000110001001110:begin data = code ^ 80'b00000000000010000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000100011110010:begin data = code ^ 80'b00000000000010000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000110001010:begin data = code ^ 80'b00000000000010000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001101111010:begin data = code ^ 80'b00000000000010000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011011010011010:begin data = code ^ 80'b00000000000010001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111110101011010:begin data = code ^ 80'b00000000000010010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110101011011010:begin data = code ^ 80'b00000000000010100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100000110111:begin data = code ^ 80'b00000000000011000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001001011000:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1001001001011011:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1001001001011101:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1001001001010001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1001001001001001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1001001001111001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1001001000011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1001001011011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1001001101011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1001000001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1001011001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1001101001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1000001001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1011001001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1101001001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0001001001011001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0001111110110100:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0000010001101110:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0011001111011010:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0101110010110010:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1000001001100010:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1011001000101111:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1101001010110101:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0001001110000001:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0001110000000100:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0000001100001110:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0011110100011010:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0100000100110010:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1011100101100010:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1100010000101111:begin data = code ^ 80'b00000000000100000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0011111010110101:begin data = code ^ 80'b00000000000100000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0100011001101100:begin data = code ^ 80'b00000000000100000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1011011111011110:begin data = code ^ 80'b00000000000100000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1101100101010111:begin data = code ^ 80'b00000000000100000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0000010001000101:begin data = code ^ 80'b00000000000100000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0011001110001100:begin data = code ^ 80'b00000000000100000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0101110000011110:begin data = code ^ 80'b00000000000100000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1000001100111010:begin data = code ^ 80'b00000000000100000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1011000010011111:begin data = code ^ 80'b00000000000100000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1101011111010101:begin data = code ^ 80'b00000000000100000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0001100101000001:begin data = code ^ 80'b00000000000100000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0000100110000100:begin data = code ^ 80'b00000000000100000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0010100000001110:begin data = code ^ 80'b00000000000100000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0110101100011010:begin data = code ^ 80'b00000000000100000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1110110100110010:begin data = code ^ 80'b00000000000100000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0110110010001111:begin data = code ^ 80'b00000000000100000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001000011000:begin data = code ^ 80'b00000000000100000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001011011011:begin data = code ^ 80'b00000000000100000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111010110000:begin data = code ^ 80'b00000000000100000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101110001011:begin data = code ^ 80'b00000000000100000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110000010000:begin data = code ^ 80'b00000000000100000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001100100110:begin data = code ^ 80'b00000000000100000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111110101001010:begin data = code ^ 80'b00000000000100000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110001111111:begin data = code ^ 80'b00000000000100000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010001111111000:begin data = code ^ 80'b00000000000100000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000100011011:begin data = code ^ 80'b00000000000100000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101010011011101:begin data = code ^ 80'b00000000000100000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001010111100:begin data = code ^ 80'b00000000000100000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001110010011:begin data = code ^ 80'b00000000000100000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000111001101:begin data = code ^ 80'b00000000000100000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001010101110001:begin data = code ^ 80'b00000000000100000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001110000001001:begin data = code ^ 80'b00000000000100000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111011111001:begin data = code ^ 80'b00000000000100000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010101100011001:begin data = code ^ 80'b00000000000100001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000011011001:begin data = code ^ 80'b00000000000100010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011101011001:begin data = code ^ 80'b00000000000100100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101010110110100:begin data = code ^ 80'b00000000000101000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110110000011:begin data = code ^ 80'b00000000000110000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100101011110:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1010100101011101:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1010100101011011:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1010100101010111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1010100101001111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1010100101111111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1010100100011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1010100111011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1010100001011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1010101101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1010110101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1010000101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1011100101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1000100101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1110100101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0010100101011111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0010010010110010:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0011111101101000:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0000100011011100:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0110011110110100:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1011100101100100:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1000100100101001:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1110100110110011:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0010100010000111:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0010011100000010:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0011100000001000:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0000011000011100:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0111101000110100:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1000001001100100:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1111111100101001:begin data = code ^ 80'b00000000001000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0000010110110011:begin data = code ^ 80'b00000000001000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0111110101101010:begin data = code ^ 80'b00000000001000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1000110011011000:begin data = code ^ 80'b00000000001000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1110001001010001:begin data = code ^ 80'b00000000001000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0011111101000011:begin data = code ^ 80'b00000000001000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0000100010001010:begin data = code ^ 80'b00000000001000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0110011100011000:begin data = code ^ 80'b00000000001000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1011100000111100:begin data = code ^ 80'b00000000001000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1000101110011001:begin data = code ^ 80'b00000000001000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1110110011010011:begin data = code ^ 80'b00000000001000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0010001001000111:begin data = code ^ 80'b00000000001000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0011001010000010:begin data = code ^ 80'b00000000001000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0001001100001000:begin data = code ^ 80'b00000000001000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000000011100:begin data = code ^ 80'b00000000001000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1101011000110100:begin data = code ^ 80'b00000000001000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0101011110001001:begin data = code ^ 80'b00000000001000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101100100011110:begin data = code ^ 80'b00000000001000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100111011101:begin data = code ^ 80'b00000000001000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110010110110110:begin data = code ^ 80'b00000000001000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000010001101:begin data = code ^ 80'b00000000001000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011100010110:begin data = code ^ 80'b00000000001000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101100000100000:begin data = code ^ 80'b00000000001000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011001001100:begin data = code ^ 80'b00000000001000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011101111001:begin data = code ^ 80'b00000000001000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100011111110:begin data = code ^ 80'b00000000001000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100101000011101:begin data = code ^ 80'b00000000001000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111111011011:begin data = code ^ 80'b00000000001000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100110111010:begin data = code ^ 80'b00000000001000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100010010101:begin data = code ^ 80'b00000000001000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010101011001011:begin data = code ^ 80'b00000000001000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111001110111:begin data = code ^ 80'b00000000001000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010011100001111:begin data = code ^ 80'b00000000001000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011010111111111:begin data = code ^ 80'b00000000001000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000000011111:begin data = code ^ 80'b00000000001000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101101111011111:begin data = code ^ 80'b00000000001000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110001011111:begin data = code ^ 80'b00000000001000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111010110010:begin data = code ^ 80'b00000000001001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011010000101:begin data = code ^ 80'b00000000001010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011101100000110:begin data = code ^ 80'b00000000001100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111101010010:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1101111101010001:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1101111101010111:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1101111101011011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1101111101000011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1101111101110011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1101111100010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1101111111010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1101111001010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1101110101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1101101101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1101011101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1100111101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1111111101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1001111101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0101111101010011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0101001010111110:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0100100101100100:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0111111011010000:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0001000110111000:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1100111101101000:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1111111100100101:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1001111110111111:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0101111010001011:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0101000100001110:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0100111000000100:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0111000000010000:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0000110000111000:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1111010001101000:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1000100100100101:begin data = code ^ 80'b00000000010000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0111001110111111:begin data = code ^ 80'b00000000010000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0000101101100110:begin data = code ^ 80'b00000000010000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1111101011010100:begin data = code ^ 80'b00000000010000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1001010001011101:begin data = code ^ 80'b00000000010000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0100100101001111:begin data = code ^ 80'b00000000010000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0111111010000110:begin data = code ^ 80'b00000000010000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0001000100010100:begin data = code ^ 80'b00000000010000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1100111000110000:begin data = code ^ 80'b00000000010000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1111110110010101:begin data = code ^ 80'b00000000010000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1001101011011111:begin data = code ^ 80'b00000000010000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0101010001001011:begin data = code ^ 80'b00000000010000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0100010010001110:begin data = code ^ 80'b00000000010000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0110010100000100:begin data = code ^ 80'b00000000010000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011000010000:begin data = code ^ 80'b00000000010000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000000111000:begin data = code ^ 80'b00000000010000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000110000101:begin data = code ^ 80'b00000000010000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111100010010:begin data = code ^ 80'b00000000010000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111111010001:begin data = code ^ 80'b00000000010000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001110111010:begin data = code ^ 80'b00000000010000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100011010000001:begin data = code ^ 80'b00000000010000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000100011010:begin data = code ^ 80'b00000000010000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111000101100:begin data = code ^ 80'b00000000010000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011000001000000:begin data = code ^ 80'b00000000010000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000000101110101:begin data = code ^ 80'b00000000010000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111011110010:begin data = code ^ 80'b00000000010000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110000010001:begin data = code ^ 80'b00000000010000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100111010111:begin data = code ^ 80'b00000000010000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111110110110:begin data = code ^ 80'b00000000010000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111010011001:begin data = code ^ 80'b00000000010000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101110011000111:begin data = code ^ 80'b00000000010000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101100001111011:begin data = code ^ 80'b00000000010000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000100000011:begin data = code ^ 80'b00000000010000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001111110011:begin data = code ^ 80'b00000000010000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110011000010011:begin data = code ^ 80'b00000000010000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010110111010011:begin data = code ^ 80'b00000000010000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011101001010011:begin data = code ^ 80'b00000000010000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100010111110:begin data = code ^ 80'b00000000010001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000010001001:begin data = code ^ 80'b00000000010010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110100001010:begin data = code ^ 80'b00000000010100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011000001100:begin data = code ^ 80'b00000000011000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001101001010:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0011001101001001:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0011001101001111:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0011001101000011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0011001101011011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0011001101101011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0011001100001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0011001111001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0011001001001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0011000101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0011011101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0011101101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0010001101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0001001101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0111001101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1011001101001011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1011111010100110:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1010010101111100:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1001001011001000:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1111110110100000:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0010001101110000:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0001001100111101:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0111001110100111:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1011001010010011:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1011110100010110:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1010001000011100:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1001110000001000:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1110000000100000:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0001100001110000:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0110010100111101:begin data = code ^ 80'b00000000100000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1001111110100111:begin data = code ^ 80'b00000000100000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1110011101111110:begin data = code ^ 80'b00000000100000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0001011011001100:begin data = code ^ 80'b00000000100000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0111100001000101:begin data = code ^ 80'b00000000100000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1010010101010111:begin data = code ^ 80'b00000000100000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1001001010011110:begin data = code ^ 80'b00000000100000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1111110100001100:begin data = code ^ 80'b00000000100000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0010001000101000:begin data = code ^ 80'b00000000100000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0001000110001101:begin data = code ^ 80'b00000000100000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0111011011000111:begin data = code ^ 80'b00000000100000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1011100001010011:begin data = code ^ 80'b00000000100000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1010100010010110:begin data = code ^ 80'b00000000100000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1000100100011100:begin data = code ^ 80'b00000000100000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1100101000001000:begin data = code ^ 80'b00000000100000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110000100000:begin data = code ^ 80'b00000000100000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110110011101:begin data = code ^ 80'b00000000100000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001100001010:begin data = code ^ 80'b00000000100000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101001111001001:begin data = code ^ 80'b00000000100000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111111110100010:begin data = code ^ 80'b00000000100000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010101010011001:begin data = code ^ 80'b00000000100000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000110100000010:begin data = code ^ 80'b00000000100000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001000110100:begin data = code ^ 80'b00000000100000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101110001011000:begin data = code ^ 80'b00000000100000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110110101101101:begin data = code ^ 80'b00000000100000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001011101010:begin data = code ^ 80'b00000000100000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000000001001:begin data = code ^ 80'b00000000100000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111010111001111:begin data = code ^ 80'b00000000100000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001110101110:begin data = code ^ 80'b00000000100000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001010000001:begin data = code ^ 80'b00000000100000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000011011111:begin data = code ^ 80'b00000000100000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011010001100011:begin data = code ^ 80'b00000000100000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011110100011011:begin data = code ^ 80'b00000000100000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111111101011:begin data = code ^ 80'b00000000100000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101000001011:begin data = code ^ 80'b00000000100000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100000111001011:begin data = code ^ 80'b00000000100000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101011001001011:begin data = code ^ 80'b00000000100000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111010010100110:begin data = code ^ 80'b00000000100001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110010010001:begin data = code ^ 80'b00000000100010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000100010010:begin data = code ^ 80'b00000000100100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001101000010100:begin data = code ^ 80'b00000000101000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110110000011000:begin data = code ^ 80'b00000000110000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011010010111:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0110011010010100:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0110011010010010:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0110011010011110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0110011010000110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0110011010110110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0110011011010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0110011000010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0110011110010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0110010010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0110001010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0110111010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0111011010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0100011010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0010011010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1110011010010110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1110101101111011:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1111000010100001:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1100011100010101:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1010100001111101:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0111011010101101:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0100011011100000:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0010011001111010:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1110011101001110:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1110100011001011:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1111011111000001:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1100100111010101:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1011010111111101:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0100110110101101:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0011000011100000:begin data = code ^ 80'b00000001000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1100101001111010:begin data = code ^ 80'b00000001000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1011001010100011:begin data = code ^ 80'b00000001000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0100001100010001:begin data = code ^ 80'b00000001000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0010110110011000:begin data = code ^ 80'b00000001000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1111000010001010:begin data = code ^ 80'b00000001000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1100011101000011:begin data = code ^ 80'b00000001000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1010100011010001:begin data = code ^ 80'b00000001000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0111011111110101:begin data = code ^ 80'b00000001000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0100010001010000:begin data = code ^ 80'b00000001000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0010001100011010:begin data = code ^ 80'b00000001000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1110110110001110:begin data = code ^ 80'b00000001000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1111110101001011:begin data = code ^ 80'b00000001000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1101110011000001:begin data = code ^ 80'b00000001000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1001111111010101:begin data = code ^ 80'b00000001000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100111111101:begin data = code ^ 80'b00000001000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100001000000:begin data = code ^ 80'b00000001000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011011010111:begin data = code ^ 80'b00000001000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011000010100:begin data = code ^ 80'b00000001000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010101001111111:begin data = code ^ 80'b00000001000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111101000100:begin data = code ^ 80'b00000001000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101100011011111:begin data = code ^ 80'b00000001000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001011111101001:begin data = code ^ 80'b00000001000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100110000101:begin data = code ^ 80'b00000001000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011100010110000:begin data = code ^ 80'b00000001000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101011100110111:begin data = code ^ 80'b00000001000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000010111010100:begin data = code ^ 80'b00000001000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000000010010:begin data = code ^ 80'b00000001000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011001110011:begin data = code ^ 80'b00000001000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011101011100:begin data = code ^ 80'b00000001000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110010100000010:begin data = code ^ 80'b00000001000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000110111110:begin data = code ^ 80'b00000001000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110100011000110:begin data = code ^ 80'b00000001000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111101000110110:begin data = code ^ 80'b00000001000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111111010110:begin data = code ^ 80'b00000001000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001010000010110:begin data = code ^ 80'b00000001000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000001110010110:begin data = code ^ 80'b00000001000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000101111011:begin data = code ^ 80'b00000001000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110100101001100:begin data = code ^ 80'b00000001000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111010011001111:begin data = code ^ 80'b00000001000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111111001001:begin data = code ^ 80'b00000001001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011100111000101:begin data = code ^ 80'b00000001010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101010111011101:begin data = code ^ 80'b00000001100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110100101101:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1100110100101110:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1100110100101000:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1100110100100100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1100110100111100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1100110100001100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1100110101101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1100110110101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1100110000101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1100111100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1100100100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1100010100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1101110100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1110110100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1000110100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0100110100101100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0100000011000001:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0101101100011011:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0110110010101111:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0000001111000111:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1101110100010111:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1110110101011010:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1000110111000000:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0100110011110100:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0100001101110001:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0101110001111011:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0110001001101111:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0001111001000111:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1110011000010111:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1001101101011010:begin data = code ^ 80'b00000010000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0110000111000000:begin data = code ^ 80'b00000010000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0001100100011001:begin data = code ^ 80'b00000010000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1110100010101011:begin data = code ^ 80'b00000010000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1000011000100010:begin data = code ^ 80'b00000010000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0101101100110000:begin data = code ^ 80'b00000010000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0110110011111001:begin data = code ^ 80'b00000010000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0000001101101011:begin data = code ^ 80'b00000010000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1101110001001111:begin data = code ^ 80'b00000010000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1110111111101010:begin data = code ^ 80'b00000010000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1000100010100000:begin data = code ^ 80'b00000010000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0100011000110100:begin data = code ^ 80'b00000010000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0101011011110001:begin data = code ^ 80'b00000010000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0111011101111011:begin data = code ^ 80'b00000010000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0011010001101111:begin data = code ^ 80'b00000010000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1011001001000111:begin data = code ^ 80'b00000010000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001111111010:begin data = code ^ 80'b00000010000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110101101101:begin data = code ^ 80'b00000010000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110110101110:begin data = code ^ 80'b00000010000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000111000101:begin data = code ^ 80'b00000010000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101010011111110:begin data = code ^ 80'b00000010000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111001101100101:begin data = code ^ 80'b00000010000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011110001010011:begin data = code ^ 80'b00000010000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010001000111111:begin data = code ^ 80'b00000010000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001100001010:begin data = code ^ 80'b00000010000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111110010001101:begin data = code ^ 80'b00000010000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111001101110:begin data = code ^ 80'b00000010000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101110101000:begin data = code ^ 80'b00000010000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110111001001:begin data = code ^ 80'b00000010000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110011100110:begin data = code ^ 80'b00000010000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111010111000:begin data = code ^ 80'b00000010000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100101000000100:begin data = code ^ 80'b00000010000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001101111100:begin data = code ^ 80'b00000010000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000110001100:begin data = code ^ 80'b00000010000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111010001101100:begin data = code ^ 80'b00000010000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111110101100:begin data = code ^ 80'b00000010000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010100000101100:begin data = code ^ 80'b00000010000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000101011000001:begin data = code ^ 80'b00000010000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001011110110:begin data = code ^ 80'b00000010000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111101110101:begin data = code ^ 80'b00000010000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110010001110011:begin data = code ^ 80'b00000010001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001001111111:begin data = code ^ 80'b00000010010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111111001100111:begin data = code ^ 80'b00000010100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010101110111010:begin data = code ^ 80'b00000011000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011110110100:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0001011110110111:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0001011110110001:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0001011110111101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0001011110100101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0001011110010101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0001011111110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0001011100110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0001011010110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0001010110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0001001110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0001111110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0000011110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0011011110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0101011110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1001011110110101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1001101001011000:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1000000110000010:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1011011000110110:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1101100101011110:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0000011110001110:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0011011111000011:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0101011101011001:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1001011001101101:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1001100111101000:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1000011011100010:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1011100011110110:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1100010011011110:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0011110010001110:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0100000111000011:begin data = code ^ 80'b00000100000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1011101101011001:begin data = code ^ 80'b00000100000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1100001110000000:begin data = code ^ 80'b00000100000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0011001000110010:begin data = code ^ 80'b00000100000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0101110010111011:begin data = code ^ 80'b00000100000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1000000110101001:begin data = code ^ 80'b00000100000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1011011001100000:begin data = code ^ 80'b00000100000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1101100111110010:begin data = code ^ 80'b00000100000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0000011011010110:begin data = code ^ 80'b00000100000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0011010101110011:begin data = code ^ 80'b00000100000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0101001000111001:begin data = code ^ 80'b00000100000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1001110010101101:begin data = code ^ 80'b00000100000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1000110001101000:begin data = code ^ 80'b00000100000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1010110111100010:begin data = code ^ 80'b00000100000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111011110110:begin data = code ^ 80'b00000100000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0110100011011110:begin data = code ^ 80'b00000100000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1110100101100011:begin data = code ^ 80'b00000100000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011111110100:begin data = code ^ 80'b00000100000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011100110111:begin data = code ^ 80'b00000100000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101101101011100:begin data = code ^ 80'b00000100000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111001100111:begin data = code ^ 80'b00000100000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100111111100:begin data = code ^ 80'b00000100000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110011011001010:begin data = code ^ 80'b00000100000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111100010100110:begin data = code ^ 80'b00000100000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100110010011:begin data = code ^ 80'b00000100000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011000010100:begin data = code ^ 80'b00000100000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111010011110111:begin data = code ^ 80'b00000100000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000100110001:begin data = code ^ 80'b00000100000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011101010000:begin data = code ^ 80'b00000100000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011001111111:begin data = code ^ 80'b00000100000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001010000100001:begin data = code ^ 80'b00000100000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000010011101:begin data = code ^ 80'b00000100000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100111100101:begin data = code ^ 80'b00000100000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000101100010101:begin data = code ^ 80'b00000100000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111011110101:begin data = code ^ 80'b00000100000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110010100110101:begin data = code ^ 80'b00000100000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111001010110101:begin data = code ^ 80'b00000100000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000001011000:begin data = code ^ 80'b00000100000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100001101111:begin data = code ^ 80'b00000100000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010111101100:begin data = code ^ 80'b00000100000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111011101010:begin data = code ^ 80'b00000100001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100011100110:begin data = code ^ 80'b00000100010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010010011111110:begin data = code ^ 80'b00000100100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000100100011:begin data = code ^ 80'b00000101000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101101010011001:begin data = code ^ 80'b00000110000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111101101011:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0010111101101000:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0010111101101110:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0010111101100010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0010111101111010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0010111101001010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0010111100101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0010111111101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0010111001101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0010110101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0010101101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0010011101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0011111101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0000111101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0110111101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1010111101101010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1010001010000111:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1011100101011101:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1000111011101001:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1110000110000001:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0011111101010001:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0000111100011100:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0110111110000110:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1010111010110010:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1010000100110111:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1011111000111101:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1000000000101001:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1111110000000001:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0000010001010001:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0111100100011100:begin data = code ^ 80'b00001000000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1000001110000110:begin data = code ^ 80'b00001000000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1111101101011111:begin data = code ^ 80'b00001000000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0000101011101101:begin data = code ^ 80'b00001000000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0110010001100100:begin data = code ^ 80'b00001000000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1011100101110110:begin data = code ^ 80'b00001000000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1000111010111111:begin data = code ^ 80'b00001000000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1110000100101101:begin data = code ^ 80'b00001000000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0011111000001001:begin data = code ^ 80'b00001000000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0000110110101100:begin data = code ^ 80'b00001000000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0110101011100110:begin data = code ^ 80'b00001000000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1010010001110010:begin data = code ^ 80'b00001000000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1011010010110111:begin data = code ^ 80'b00001000000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1001010100111101:begin data = code ^ 80'b00001000000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1101011000101001:begin data = code ^ 80'b00001000000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000000000001:begin data = code ^ 80'b00001000000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000110111100:begin data = code ^ 80'b00001000000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111100101011:begin data = code ^ 80'b00001000000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111111101000:begin data = code ^ 80'b00001000000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001110000011:begin data = code ^ 80'b00001000000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011011010111000:begin data = code ^ 80'b00001000000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000100100011:begin data = code ^ 80'b00001000000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111000010101:begin data = code ^ 80'b00001000000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100000001111001:begin data = code ^ 80'b00001000000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000101001100:begin data = code ^ 80'b00001000000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001111011001011:begin data = code ^ 80'b00001000000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110000101000:begin data = code ^ 80'b00001000000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110100111101110:begin data = code ^ 80'b00001000000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111110001111:begin data = code ^ 80'b00001000000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111010100000:begin data = code ^ 80'b00001000000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110011111110:begin data = code ^ 80'b00001000000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010100001000010:begin data = code ^ 80'b00001000000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000100111010:begin data = code ^ 80'b00001000000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001111001010:begin data = code ^ 80'b00001000000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011000101010:begin data = code ^ 80'b00001000000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101110111101010:begin data = code ^ 80'b00001000000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100101001101010:begin data = code ^ 80'b00001000000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110100010000111:begin data = code ^ 80'b00001000000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000010110000:begin data = code ^ 80'b00001000000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110100110011:begin data = code ^ 80'b00001000000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011000110101:begin data = code ^ 80'b00001000001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000000111001:begin data = code ^ 80'b00001000010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001110000100001:begin data = code ^ 80'b00001000100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100111111100:begin data = code ^ 80'b00001001000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001001000110:begin data = code ^ 80'b00001010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100011011111:begin data = code ^ 80'b00001100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111011010101:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0101111011010110:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0101111011010000:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0101111011011100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0101111011000100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0101111011110100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0101111010010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0101111001010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0101111111010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0101110011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0101101011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0101011011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0100111011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0111111011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0001111011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1101111011010100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1101001100111001:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1100100011100011:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1111111101010111:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1001000000111111:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0100111011101111:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0111111010100010:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0001111000111000:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1101111100001100:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1101000010001001:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1100111110000011:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1111000110010111:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1000110110111111:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0111010111101111:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0000100010100010:begin data = code ^ 80'b00010000000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1111001000111000:begin data = code ^ 80'b00010000000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1000101011100001:begin data = code ^ 80'b00010000000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0111101101010011:begin data = code ^ 80'b00010000000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0001010111011010:begin data = code ^ 80'b00010000000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1100100011001000:begin data = code ^ 80'b00010000000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1111111100000001:begin data = code ^ 80'b00010000000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1001000010010011:begin data = code ^ 80'b00010000000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0100111110110111:begin data = code ^ 80'b00010000000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0111110000010010:begin data = code ^ 80'b00010000000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0001101101011000:begin data = code ^ 80'b00010000000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1101010111001100:begin data = code ^ 80'b00010000000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1100010100001001:begin data = code ^ 80'b00010000000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1110010010000011:begin data = code ^ 80'b00010000000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1010011110010111:begin data = code ^ 80'b00010000000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0010000110111111:begin data = code ^ 80'b00010000000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000000000010:begin data = code ^ 80'b00010000000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111010010101:begin data = code ^ 80'b00010000000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111001010110:begin data = code ^ 80'b00010000000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001000111101:begin data = code ^ 80'b00010000000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011100000110:begin data = code ^ 80'b00010000000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000010011101:begin data = code ^ 80'b00010000000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010111110101011:begin data = code ^ 80'b00010000000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000111000111:begin data = code ^ 80'b00010000000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000011110010:begin data = code ^ 80'b00010000000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111101110101:begin data = code ^ 80'b00010000000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011110110010110:begin data = code ^ 80'b00010000000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100001010000:begin data = code ^ 80'b00010000000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111000110001:begin data = code ^ 80'b00010000000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111100011110:begin data = code ^ 80'b00010000000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101110101000000:begin data = code ^ 80'b00010000000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101100111111100:begin data = code ^ 80'b00010000000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000010000100:begin data = code ^ 80'b00010000000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001001110100:begin data = code ^ 80'b00010000000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011110010100:begin data = code ^ 80'b00010000000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110001010100:begin data = code ^ 80'b00010000000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011101111010100:begin data = code ^ 80'b00010000000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001100100111001:begin data = code ^ 80'b00010000000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101000100001110:begin data = code ^ 80'b00010000000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110010001101:begin data = code ^ 80'b00010000000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011110001011:begin data = code ^ 80'b00010000001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000110000111:begin data = code ^ 80'b00010000010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110110110011111:begin data = code ^ 80'b00010000100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011100001000010:begin data = code ^ 80'b00010001000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001111111000:begin data = code ^ 80'b00010010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100101100001:begin data = code ^ 80'b00010100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000110111110:begin data = code ^ 80'b00011000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110110101001:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1011110110101010:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1011110110101100:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1011110110100000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1011110110111000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1011110110001000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1011110111101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1011110100101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1011110010101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1011111110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1011100110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1011010110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1010110110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1001110110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1111110110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0011110110101000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0011000001000101:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0010101110011111:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0001110000101011:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0111001101000011:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1010110110010011:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1001110111011110:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1111110101000100:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0011110001110000:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0011001111110101:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0010110011111111:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0001001011101011:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0110111011000011:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1001011010010011:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1110101111011110:begin data = code ^ 80'b00100000000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0001000101000100:begin data = code ^ 80'b00100000000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0110100110011101:begin data = code ^ 80'b00100000000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1001100000101111:begin data = code ^ 80'b00100000000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1111011010100110:begin data = code ^ 80'b00100000000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0010101110110100:begin data = code ^ 80'b00100000000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0001110001111101:begin data = code ^ 80'b00100000000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0111001111101111:begin data = code ^ 80'b00100000000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1010110011001011:begin data = code ^ 80'b00100000000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1001111101101110:begin data = code ^ 80'b00100000000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1111100000100100:begin data = code ^ 80'b00100000000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0011011010110000:begin data = code ^ 80'b00100000000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0010011001110101:begin data = code ^ 80'b00100000000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0000011111111111:begin data = code ^ 80'b00100000000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0100010011101011:begin data = code ^ 80'b00100000000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1100001011000011:begin data = code ^ 80'b00100000000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0100001101111110:begin data = code ^ 80'b00100000000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100110111101001:begin data = code ^ 80'b00100000000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101110100101010:begin data = code ^ 80'b00100000000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000101000001:begin data = code ^ 80'b00100000000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010010001111010:begin data = code ^ 80'b00100000000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001111100001:begin data = code ^ 80'b00100000000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100110011010111:begin data = code ^ 80'b00100000000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101001010111011:begin data = code ^ 80'b00100000000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001110001110:begin data = code ^ 80'b00100000000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000110000001001:begin data = code ^ 80'b00100000000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111011101010:begin data = code ^ 80'b00100000000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111101100101100:begin data = code ^ 80'b00100000000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110101001101:begin data = code ^ 80'b00100000000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011110001100010:begin data = code ^ 80'b00100000000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111000111100:begin data = code ^ 80'b00100000000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011101010000000:begin data = code ^ 80'b00100000000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011001111111000:begin data = code ^ 80'b00100000000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010000100001000:begin data = code ^ 80'b00100000000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010011101000:begin data = code ^ 80'b00100000000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111100101000:begin data = code ^ 80'b00100000000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101100010101000:begin data = code ^ 80'b00100000000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111101001000101:begin data = code ^ 80'b00100000000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011001001110010:begin data = code ^ 80'b00100000000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010111111110001:begin data = code ^ 80'b00100000000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001010011110111:begin data = code ^ 80'b00100000001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001011111011:begin data = code ^ 80'b00100000010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000111011100011:begin data = code ^ 80'b00100000100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101101100111110:begin data = code ^ 80'b00100001000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111000010000100:begin data = code ^ 80'b00100010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010101000011101:begin data = code ^ 80'b00100100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001001011000010:begin data = code ^ 80'b00101000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110001101111100:begin data = code ^ 80'b00110000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011010111100:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b1111011010111111:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b1111011010111001:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b1111011010110101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b1111011010101101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b1111011010011101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b1111011011111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b1111011000111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b1111011110111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b1111010010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b1111001010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b1111111010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b1110011010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b1101011010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b1011011010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b0111011010111101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b0111101101010000:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b0110000010001010:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b0101011100111110:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b0011100001010110:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b1110011010000110:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b1101011011001011:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b1011011001010001:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b0111011101100101:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b0111100011100000:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b0110011111101010:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b0101100111111110:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b0010010111010110:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b1101110110000110:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b1010000011001011:begin data = code ^ 80'b01000000000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b0101101001010001:begin data = code ^ 80'b01000000000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b0010001010001000:begin data = code ^ 80'b01000000000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b1101001100111010:begin data = code ^ 80'b01000000000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b1011110110110011:begin data = code ^ 80'b01000000000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b0110000010100001:begin data = code ^ 80'b01000000000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b0101011101101000:begin data = code ^ 80'b01000000000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b0011100011111010:begin data = code ^ 80'b01000000000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b1110011111011110:begin data = code ^ 80'b01000000000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b1101010001111011:begin data = code ^ 80'b01000000000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b1011001100110001:begin data = code ^ 80'b01000000000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b0111110110100101:begin data = code ^ 80'b01000000000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b0110110101100000:begin data = code ^ 80'b01000000000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b0100110011101010:begin data = code ^ 80'b01000000000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111111111110:begin data = code ^ 80'b01000000000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b1000100111010110:begin data = code ^ 80'b01000000000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b0000100001101011:begin data = code ^ 80'b01000000000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000011011111100:begin data = code ^ 80'b01000000000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001011000111111:begin data = code ^ 80'b01000000000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011101001010100:begin data = code ^ 80'b01000000000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111101101111:begin data = code ^ 80'b01000000000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100100011110100:begin data = code ^ 80'b01000000000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011111000010:begin data = code ^ 80'b01000000000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100110101110:begin data = code ^ 80'b01000000000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010100010011011:begin data = code ^ 80'b01000000000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100011100011100:begin data = code ^ 80'b01000000000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001010111111111:begin data = code ^ 80'b01000000000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011000000111001:begin data = code ^ 80'b01000000000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011001011000:begin data = code ^ 80'b01000000000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111011101110111:begin data = code ^ 80'b01000000000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111010100101001:begin data = code ^ 80'b01000000000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111000110010101:begin data = code ^ 80'b01000000000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100011101101:begin data = code ^ 80'b01000000000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110101000011101:begin data = code ^ 80'b01000000000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100111111111101:begin data = code ^ 80'b01000000000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010000111101:begin data = code ^ 80'b01000000000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001110111101:begin data = code ^ 80'b01000000000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011000101010000:begin data = code ^ 80'b01000000000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111100101100111:begin data = code ^ 80'b01000000000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110010011100100:begin data = code ^ 80'b01000000000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101111111100010:begin data = code ^ 80'b01000000001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010100111101110:begin data = code ^ 80'b01000000010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100010111110110:begin data = code ^ 80'b01000000100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000000101011:begin data = code ^ 80'b01000001000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011101110010001:begin data = code ^ 80'b01000010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110000100001000:begin data = code ^ 80'b01000100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101100111010111:begin data = code ^ 80'b01001000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010100001101001:begin data = code ^ 80'b01010000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100101100010101:begin data = code ^ 80'b01100000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000010010110:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000000001; ec = 1; end
        16'b0110000010010101:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000000010; ec = 1; end
        16'b0110000010010011:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000000100; ec = 1; end
        16'b0110000010011111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000001000; ec = 1; end
        16'b0110000010000111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000010000; ec = 1; end
        16'b0110000010110111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000000100000; ec = 1; end
        16'b0110000011010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000001000000; ec = 1; end
        16'b0110000000010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000010000000; ec = 1; end
        16'b0110000110010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000000100000000; ec = 1; end
        16'b0110001010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000001000000000; ec = 1; end
        16'b0110010010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000010000000000; ec = 1; end
        16'b0110100010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000000100000000000; ec = 1; end
        16'b0111000010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000001000000000000; ec = 1; end
        16'b0100000010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000010000000000000; ec = 1; end
        16'b0010000010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000000100000000000000; ec = 1; end
        16'b1110000010010111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000001000000000000000; ec = 1; end
        16'b1110110101111010:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000010000000000000000; ec = 1; end
        16'b1111011010100000:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000000100000000000000000; ec = 1; end
        16'b1100000100010100:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000001000000000000000000; ec = 1; end
        16'b1010111001111100:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000010000000000000000000; ec = 1; end
        16'b0111000010101100:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000000100000000000000000000; ec = 1; end
        16'b0100000011100001:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000001000000000000000000000; ec = 1; end
        16'b0010000001111011:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000010000000000000000000000; ec = 1; end
        16'b1110000101001111:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000000100000000000000000000000; ec = 1; end
        16'b1110111011001010:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000001000000000000000000000000; ec = 1; end
        16'b1111000111000000:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000010000000000000000000000000; ec = 1; end
        16'b1100111111010100:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000000100000000000000000000000000; ec = 1; end
        16'b1011001111111100:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000001000000000000000000000000000; ec = 1; end
        16'b0100101110101100:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000010000000000000000000000000000; ec = 1; end
        16'b0011011011100001:begin data = code ^ 80'b10000000000000000000000000000000000000000000000000100000000000000000000000000000; ec = 1; end
        16'b1100110001111011:begin data = code ^ 80'b10000000000000000000000000000000000000000000000001000000000000000000000000000000; ec = 1; end
        16'b1011010010100010:begin data = code ^ 80'b10000000000000000000000000000000000000000000000010000000000000000000000000000000; ec = 1; end
        16'b0100010100010000:begin data = code ^ 80'b10000000000000000000000000000000000000000000000100000000000000000000000000000000; ec = 1; end
        16'b0010101110011001:begin data = code ^ 80'b10000000000000000000000000000000000000000000001000000000000000000000000000000000; ec = 1; end
        16'b1111011010001011:begin data = code ^ 80'b10000000000000000000000000000000000000000000010000000000000000000000000000000000; ec = 1; end
        16'b1100000101000010:begin data = code ^ 80'b10000000000000000000000000000000000000000000100000000000000000000000000000000000; ec = 1; end
        16'b1010111011010000:begin data = code ^ 80'b10000000000000000000000000000000000000000001000000000000000000000000000000000000; ec = 1; end
        16'b0111000111110100:begin data = code ^ 80'b10000000000000000000000000000000000000000010000000000000000000000000000000000000; ec = 1; end
        16'b0100001001010001:begin data = code ^ 80'b10000000000000000000000000000000000000000100000000000000000000000000000000000000; ec = 1; end
        16'b0010010100011011:begin data = code ^ 80'b10000000000000000000000000000000000000001000000000000000000000000000000000000000; ec = 1; end
        16'b1110101110001111:begin data = code ^ 80'b10000000000000000000000000000000000000010000000000000000000000000000000000000000; ec = 1; end
        16'b1111101101001010:begin data = code ^ 80'b10000000000000000000000000000000000000100000000000000000000000000000000000000000; ec = 1; end
        16'b1101101011000000:begin data = code ^ 80'b10000000000000000000000000000000000001000000000000000000000000000000000000000000; ec = 1; end
        16'b1001100111010100:begin data = code ^ 80'b10000000000000000000000000000000000010000000000000000000000000000000000000000000; ec = 1; end
        16'b0001111111111100:begin data = code ^ 80'b10000000000000000000000000000000000100000000000000000000000000000000000000000000; ec = 1; end
        16'b1001111001000001:begin data = code ^ 80'b10000000000000000000000000000000001000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001000011010110:begin data = code ^ 80'b10000000000000000000000000000000010000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000000000010101:begin data = code ^ 80'b10000000000000000000000000000000100000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010110001111110:begin data = code ^ 80'b10000000000000000000000000000001000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111100101000101:begin data = code ^ 80'b10000000000000000000000000000010000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101111011011110:begin data = code ^ 80'b10000000000000000000000000000100000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001000111101000:begin data = code ^ 80'b10000000000000000000000000001000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000111110000100:begin data = code ^ 80'b10000000000000000000000000010000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111010110001:begin data = code ^ 80'b10000000000000000000000000100000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101000100110110:begin data = code ^ 80'b10000000000000000000000001000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000001111010101:begin data = code ^ 80'b10000000000000000000000010000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010011000010011:begin data = code ^ 80'b10000000000000000000000100000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000001110010:begin data = code ^ 80'b10000000000000000000001000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110000101011101:begin data = code ^ 80'b10000000000000000000010000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110001100000011:begin data = code ^ 80'b10000000000000000000100000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110011110111111:begin data = code ^ 80'b10000000000000000001000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0110111011000111:begin data = code ^ 80'b10000000000000000010000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111110000110111:begin data = code ^ 80'b10000000000000000100000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101100111010111:begin data = code ^ 80'b10000000000000001000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0001001000010111:begin data = code ^ 80'b10000000000000010000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1000010110010111:begin data = code ^ 80'b10000000000000100000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0010011101111010:begin data = code ^ 80'b10000000000001000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1110111101001101:begin data = code ^ 80'b10000000000010000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1111001011001110:begin data = code ^ 80'b10000000000100000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1100100111001000:begin data = code ^ 80'b10000000001000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1011111111000100:begin data = code ^ 80'b10000000010000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0101001111011100:begin data = code ^ 80'b10000000100000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0000011000000001:begin data = code ^ 80'b10000001000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1010110110111011:begin data = code ^ 80'b10000010000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0111011100100010:begin data = code ^ 80'b10000100000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0100111111111101:begin data = code ^ 80'b10001000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b0011111001000011:begin data = code ^ 80'b10010000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1101110100111111:begin data = code ^ 80'b10100000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        16'b1001011000101010:begin data = code ^ 80'b11000000000000000000000000000000000000000000000000000000000000000000000000000000; ec = 1; end
        default : ec = 0;
    endcase
    
    dataout = data[79 -: 64];
    
end

endmodule

module add(input [7:0] add_a,add_b,
			output [7:0] sum);

assign sum = add_a + add_b;

endmodule